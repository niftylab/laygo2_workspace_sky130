magic
tech sky130A
timestamp 1679561063
<< checkpaint >>
rect -650 -660 4106 1668
<< metal1 >>
rect 1641 844 1671 1028
rect 1785 844 1815 1028
rect 1641 -20 1671 164
rect 1785 -20 1815 164
<< metal2 >>
rect -20 978 3476 1038
rect 1656 777 1800 807
rect 2289 417 2535 447
rect 1656 201 1800 231
rect -20 -30 3476 30
<< metal3 >>
rect 57 201 87 648
rect 129 417 159 807
rect 417 360 447 648
rect 777 417 807 663
rect 1425 417 1455 807
rect 2217 417 2247 663
rect 633 201 663 375
rect 2001 201 2031 375
rect 2289 129 2319 447
rect 2505 345 2535 447
rect 3297 216 3327 792
<< metal4 >>
rect 129 417 807 447
rect 1425 417 2247 447
rect 57 201 2031 231
use logic_generated_inv_2x  inv0 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 0 0 1 0
box -20 -30 308 1038
use logic_generated_inv_12x  inv1 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 2448 0 1 0
box -20 -30 1028 1038
use logic_generated_latch_2ck_2x  latch0 magic_layout/logic_generated
timestamp 1679560976
transform 1 0 288 0 1 0
box -20 -30 1316 1038
use ntap_fast_boundary  MNT0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825115
transform 1 0 1584 0 1 0
box 0 0 72 512
use ntap_fast_boundary  MNT0_IBNDR0
timestamp 1655825115
transform 1 0 1800 0 1 0
box 0 0 72 512
use ntap_fast_center_nf2_v2  MNT0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656694979
transform 1 0 1656 0 1 0
box -36 143 180 342
use via_M1_M2_0  MNT0_IVTAP10 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1728 0 1 216
box -16 -16 16 16
use via_M1_M2_1  MNT0_IVTIETAP10 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 1656 0 1 0
box -16 -16 16 16
use ptap_fast_boundary  MPT0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825477
transform 1 0 1584 0 -1 1008
box 0 0 84 512
use ptap_fast_boundary  MPT0_IBNDR0
timestamp 1655825477
transform 1 0 1800 0 -1 1008
box 0 0 84 512
use ptap_fast_center_nf2_v2  MPT0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656699071
transform 1 0 1656 0 -1 1008
box -36 66 180 342
use via_M1_M2_0  MPT0_IVTAP10
timestamp 1647525606
transform 1 0 1728 0 -1 792
box -16 -16 16 16
use via_M1_M2_1  MPT0_IVTIETAP10
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 1656 0 -1 1008
box -16 -16 16 16
use logic_generated_nand_2x  nand0 magic_layout/logic_generated
timestamp 1679560872
transform 1 0 1872 0 1 0
box -20 -30 596 1038
use via_M3_M4_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 72 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_3
timestamp 1647526059
transform 1 0 648 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_5
timestamp 1647526059
transform 1 0 2016 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_8
timestamp 1647526059
transform 1 0 144 0 1 432
box -19 -19 19 19
use via_M3_M4_0  NoName_10
timestamp 1647526059
transform 1 0 792 0 1 432
box -19 -19 19 19
use via_M3_M4_0  NoName_13
timestamp 1647526059
transform 1 0 1440 0 1 432
box -19 -19 19 19
use via_M3_M4_0  NoName_15
timestamp 1647526059
transform 1 0 2232 0 1 432
box -19 -19 19 19
use via_M2_M3_0  NoName_18 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 2304 0 1 432
box -19 -19 19 19
use via_M2_M3_0  NoName_20
timestamp 1647525786
transform 1 0 2520 0 1 432
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 CK_I
port 1 nsew
flabel metal3 3312 504 3312 504 0 FreeSans 240 90 0 0 CK_O
port 2 nsew
flabel metal3 432 504 432 504 0 FreeSans 240 90 0 0 EN
port 3 nsew
flabel metal2 1728 1008 1728 1008 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel metal2 1728 0 1728 0 0 FreeSans 480 0 0 0 VSS
port 5 nsew
<< end >>
