magic
tech sky130A
magscale 1 2
timestamp 1655978049
<< nwell >>
rect 0 1332 6336 1884
<< pwell >>
rect 0 372 6336 684
<< pmos >>
rect 200 1368 230 1848
rect 344 1368 374 1848
rect 776 1368 806 1848
rect 920 1368 950 1848
rect 1352 1368 1382 1848
rect 1496 1368 1526 1848
rect 1928 1368 1958 1848
rect 2072 1368 2102 1848
rect 2504 1368 2534 1848
rect 2648 1368 2678 1848
rect 3368 1368 3398 1848
rect 3512 1368 3542 1848
rect 3944 1368 3974 1848
rect 4088 1368 4118 1848
rect 4520 1368 4550 1848
rect 4664 1368 4694 1848
rect 5096 1368 5126 1848
rect 5240 1368 5270 1848
rect 5960 1368 5990 1848
rect 6104 1368 6134 1848
<< nmoslvt >>
rect 200 408 230 648
rect 344 408 374 648
rect 776 408 806 648
rect 920 408 950 648
rect 1352 408 1382 648
rect 1496 408 1526 648
rect 1928 408 1958 648
rect 2072 408 2102 648
rect 2504 408 2534 648
rect 2648 408 2678 648
rect 3368 408 3398 648
rect 3512 408 3542 648
rect 3944 408 3974 648
rect 4088 408 4118 648
rect 4520 408 4550 648
rect 4664 408 4694 648
rect 5096 408 5126 648
rect 5240 408 5270 648
rect 5960 408 5990 648
rect 6104 408 6134 648
<< ndiff >>
rect 88 598 200 648
rect 88 558 124 598
rect 164 558 200 598
rect 88 498 200 558
rect 88 458 124 498
rect 164 458 200 498
rect 88 408 200 458
rect 230 598 344 648
rect 230 558 268 598
rect 308 558 344 598
rect 230 498 344 558
rect 230 458 268 498
rect 308 458 344 498
rect 230 408 344 458
rect 374 598 488 648
rect 374 558 412 598
rect 452 558 488 598
rect 374 498 488 558
rect 374 458 412 498
rect 452 458 488 498
rect 374 408 488 458
rect 664 598 776 648
rect 664 558 700 598
rect 740 558 776 598
rect 664 498 776 558
rect 664 458 700 498
rect 740 458 776 498
rect 664 408 776 458
rect 806 598 920 648
rect 806 558 844 598
rect 884 558 920 598
rect 806 498 920 558
rect 806 458 844 498
rect 884 458 920 498
rect 806 408 920 458
rect 950 598 1064 648
rect 950 558 988 598
rect 1028 558 1064 598
rect 950 498 1064 558
rect 950 458 988 498
rect 1028 458 1064 498
rect 950 408 1064 458
rect 1240 598 1352 648
rect 1240 558 1276 598
rect 1316 558 1352 598
rect 1240 498 1352 558
rect 1240 458 1276 498
rect 1316 458 1352 498
rect 1240 408 1352 458
rect 1382 598 1496 648
rect 1382 558 1420 598
rect 1460 558 1496 598
rect 1382 498 1496 558
rect 1382 458 1420 498
rect 1460 458 1496 498
rect 1382 408 1496 458
rect 1526 598 1640 648
rect 1526 558 1564 598
rect 1604 558 1640 598
rect 1526 498 1640 558
rect 1526 458 1564 498
rect 1604 458 1640 498
rect 1526 408 1640 458
rect 1816 598 1928 648
rect 1816 558 1852 598
rect 1892 558 1928 598
rect 1816 498 1928 558
rect 1816 458 1852 498
rect 1892 458 1928 498
rect 1816 408 1928 458
rect 1958 598 2072 648
rect 1958 558 1996 598
rect 2036 558 2072 598
rect 1958 498 2072 558
rect 1958 458 1996 498
rect 2036 458 2072 498
rect 1958 408 2072 458
rect 2102 598 2216 648
rect 2102 558 2140 598
rect 2180 558 2216 598
rect 2102 498 2216 558
rect 2102 458 2140 498
rect 2180 458 2216 498
rect 2102 408 2216 458
rect 2392 598 2504 648
rect 2392 558 2428 598
rect 2468 558 2504 598
rect 2392 498 2504 558
rect 2392 458 2428 498
rect 2468 458 2504 498
rect 2392 408 2504 458
rect 2534 598 2648 648
rect 2534 558 2572 598
rect 2612 558 2648 598
rect 2534 498 2648 558
rect 2534 458 2572 498
rect 2612 458 2648 498
rect 2534 408 2648 458
rect 2678 598 2792 648
rect 2678 558 2716 598
rect 2756 558 2792 598
rect 2678 498 2792 558
rect 2678 458 2716 498
rect 2756 458 2792 498
rect 2678 408 2792 458
rect 3256 598 3368 648
rect 3256 558 3292 598
rect 3332 558 3368 598
rect 3256 498 3368 558
rect 3256 458 3292 498
rect 3332 458 3368 498
rect 3256 408 3368 458
rect 3398 598 3512 648
rect 3398 558 3436 598
rect 3476 558 3512 598
rect 3398 498 3512 558
rect 3398 458 3436 498
rect 3476 458 3512 498
rect 3398 408 3512 458
rect 3542 598 3656 648
rect 3542 558 3580 598
rect 3620 558 3656 598
rect 3542 498 3656 558
rect 3542 458 3580 498
rect 3620 458 3656 498
rect 3542 408 3656 458
rect 3832 598 3944 648
rect 3832 558 3868 598
rect 3908 558 3944 598
rect 3832 498 3944 558
rect 3832 458 3868 498
rect 3908 458 3944 498
rect 3832 408 3944 458
rect 3974 598 4088 648
rect 3974 558 4012 598
rect 4052 558 4088 598
rect 3974 498 4088 558
rect 3974 458 4012 498
rect 4052 458 4088 498
rect 3974 408 4088 458
rect 4118 598 4232 648
rect 4118 558 4156 598
rect 4196 558 4232 598
rect 4118 498 4232 558
rect 4118 458 4156 498
rect 4196 458 4232 498
rect 4118 408 4232 458
rect 4408 598 4520 648
rect 4408 558 4444 598
rect 4484 558 4520 598
rect 4408 498 4520 558
rect 4408 458 4444 498
rect 4484 458 4520 498
rect 4408 408 4520 458
rect 4550 598 4664 648
rect 4550 558 4588 598
rect 4628 558 4664 598
rect 4550 498 4664 558
rect 4550 458 4588 498
rect 4628 458 4664 498
rect 4550 408 4664 458
rect 4694 598 4808 648
rect 4694 558 4732 598
rect 4772 558 4808 598
rect 4694 498 4808 558
rect 4694 458 4732 498
rect 4772 458 4808 498
rect 4694 408 4808 458
rect 4984 598 5096 648
rect 4984 558 5020 598
rect 5060 558 5096 598
rect 4984 498 5096 558
rect 4984 458 5020 498
rect 5060 458 5096 498
rect 4984 408 5096 458
rect 5126 598 5240 648
rect 5126 558 5164 598
rect 5204 558 5240 598
rect 5126 498 5240 558
rect 5126 458 5164 498
rect 5204 458 5240 498
rect 5126 408 5240 458
rect 5270 598 5384 648
rect 5270 558 5308 598
rect 5348 558 5384 598
rect 5270 498 5384 558
rect 5270 458 5308 498
rect 5348 458 5384 498
rect 5270 408 5384 458
rect 5848 598 5960 648
rect 5848 558 5884 598
rect 5924 558 5960 598
rect 5848 498 5960 558
rect 5848 458 5884 498
rect 5924 458 5960 498
rect 5848 408 5960 458
rect 5990 598 6104 648
rect 5990 558 6028 598
rect 6068 558 6104 598
rect 5990 498 6104 558
rect 5990 458 6028 498
rect 6068 458 6104 498
rect 5990 408 6104 458
rect 6134 598 6248 648
rect 6134 558 6172 598
rect 6212 558 6248 598
rect 6134 498 6248 558
rect 6134 458 6172 498
rect 6212 458 6248 498
rect 6134 408 6248 458
<< pdiff >>
rect 88 1778 200 1848
rect 88 1738 124 1778
rect 164 1738 200 1778
rect 88 1678 200 1738
rect 88 1638 124 1678
rect 164 1638 200 1678
rect 88 1578 200 1638
rect 88 1538 124 1578
rect 164 1538 200 1578
rect 88 1478 200 1538
rect 88 1438 124 1478
rect 164 1438 200 1478
rect 88 1368 200 1438
rect 230 1778 344 1848
rect 230 1738 268 1778
rect 308 1738 344 1778
rect 230 1678 344 1738
rect 230 1638 268 1678
rect 308 1638 344 1678
rect 230 1578 344 1638
rect 230 1538 268 1578
rect 308 1538 344 1578
rect 230 1478 344 1538
rect 230 1438 268 1478
rect 308 1438 344 1478
rect 230 1368 344 1438
rect 374 1778 488 1848
rect 374 1738 412 1778
rect 452 1738 488 1778
rect 374 1678 488 1738
rect 374 1638 412 1678
rect 452 1638 488 1678
rect 374 1578 488 1638
rect 374 1538 412 1578
rect 452 1538 488 1578
rect 374 1478 488 1538
rect 374 1438 412 1478
rect 452 1438 488 1478
rect 374 1368 488 1438
rect 664 1778 776 1848
rect 664 1738 700 1778
rect 740 1738 776 1778
rect 664 1678 776 1738
rect 664 1638 700 1678
rect 740 1638 776 1678
rect 664 1578 776 1638
rect 664 1538 700 1578
rect 740 1538 776 1578
rect 664 1478 776 1538
rect 664 1438 700 1478
rect 740 1438 776 1478
rect 664 1368 776 1438
rect 806 1778 920 1848
rect 806 1738 844 1778
rect 884 1738 920 1778
rect 806 1678 920 1738
rect 806 1638 844 1678
rect 884 1638 920 1678
rect 806 1578 920 1638
rect 806 1538 844 1578
rect 884 1538 920 1578
rect 806 1478 920 1538
rect 806 1438 844 1478
rect 884 1438 920 1478
rect 806 1368 920 1438
rect 950 1778 1064 1848
rect 950 1738 988 1778
rect 1028 1738 1064 1778
rect 950 1678 1064 1738
rect 950 1638 988 1678
rect 1028 1638 1064 1678
rect 950 1578 1064 1638
rect 950 1538 988 1578
rect 1028 1538 1064 1578
rect 950 1478 1064 1538
rect 950 1438 988 1478
rect 1028 1438 1064 1478
rect 950 1368 1064 1438
rect 1240 1778 1352 1848
rect 1240 1738 1276 1778
rect 1316 1738 1352 1778
rect 1240 1678 1352 1738
rect 1240 1638 1276 1678
rect 1316 1638 1352 1678
rect 1240 1578 1352 1638
rect 1240 1538 1276 1578
rect 1316 1538 1352 1578
rect 1240 1478 1352 1538
rect 1240 1438 1276 1478
rect 1316 1438 1352 1478
rect 1240 1368 1352 1438
rect 1382 1778 1496 1848
rect 1382 1738 1420 1778
rect 1460 1738 1496 1778
rect 1382 1678 1496 1738
rect 1382 1638 1420 1678
rect 1460 1638 1496 1678
rect 1382 1578 1496 1638
rect 1382 1538 1420 1578
rect 1460 1538 1496 1578
rect 1382 1478 1496 1538
rect 1382 1438 1420 1478
rect 1460 1438 1496 1478
rect 1382 1368 1496 1438
rect 1526 1778 1640 1848
rect 1526 1738 1564 1778
rect 1604 1738 1640 1778
rect 1526 1678 1640 1738
rect 1526 1638 1564 1678
rect 1604 1638 1640 1678
rect 1526 1578 1640 1638
rect 1526 1538 1564 1578
rect 1604 1538 1640 1578
rect 1526 1478 1640 1538
rect 1526 1438 1564 1478
rect 1604 1438 1640 1478
rect 1526 1368 1640 1438
rect 1816 1778 1928 1848
rect 1816 1738 1852 1778
rect 1892 1738 1928 1778
rect 1816 1678 1928 1738
rect 1816 1638 1852 1678
rect 1892 1638 1928 1678
rect 1816 1578 1928 1638
rect 1816 1538 1852 1578
rect 1892 1538 1928 1578
rect 1816 1478 1928 1538
rect 1816 1438 1852 1478
rect 1892 1438 1928 1478
rect 1816 1368 1928 1438
rect 1958 1778 2072 1848
rect 1958 1738 1996 1778
rect 2036 1738 2072 1778
rect 1958 1678 2072 1738
rect 1958 1638 1996 1678
rect 2036 1638 2072 1678
rect 1958 1578 2072 1638
rect 1958 1538 1996 1578
rect 2036 1538 2072 1578
rect 1958 1478 2072 1538
rect 1958 1438 1996 1478
rect 2036 1438 2072 1478
rect 1958 1368 2072 1438
rect 2102 1778 2216 1848
rect 2102 1738 2140 1778
rect 2180 1738 2216 1778
rect 2102 1678 2216 1738
rect 2102 1638 2140 1678
rect 2180 1638 2216 1678
rect 2102 1578 2216 1638
rect 2102 1538 2140 1578
rect 2180 1538 2216 1578
rect 2102 1478 2216 1538
rect 2102 1438 2140 1478
rect 2180 1438 2216 1478
rect 2102 1368 2216 1438
rect 2392 1778 2504 1848
rect 2392 1738 2428 1778
rect 2468 1738 2504 1778
rect 2392 1678 2504 1738
rect 2392 1638 2428 1678
rect 2468 1638 2504 1678
rect 2392 1578 2504 1638
rect 2392 1538 2428 1578
rect 2468 1538 2504 1578
rect 2392 1478 2504 1538
rect 2392 1438 2428 1478
rect 2468 1438 2504 1478
rect 2392 1368 2504 1438
rect 2534 1778 2648 1848
rect 2534 1738 2572 1778
rect 2612 1738 2648 1778
rect 2534 1678 2648 1738
rect 2534 1638 2572 1678
rect 2612 1638 2648 1678
rect 2534 1578 2648 1638
rect 2534 1538 2572 1578
rect 2612 1538 2648 1578
rect 2534 1478 2648 1538
rect 2534 1438 2572 1478
rect 2612 1438 2648 1478
rect 2534 1368 2648 1438
rect 2678 1778 2792 1848
rect 2678 1738 2716 1778
rect 2756 1738 2792 1778
rect 2678 1678 2792 1738
rect 2678 1638 2716 1678
rect 2756 1638 2792 1678
rect 2678 1578 2792 1638
rect 2678 1538 2716 1578
rect 2756 1538 2792 1578
rect 2678 1478 2792 1538
rect 2678 1438 2716 1478
rect 2756 1438 2792 1478
rect 2678 1368 2792 1438
rect 3256 1778 3368 1848
rect 3256 1738 3292 1778
rect 3332 1738 3368 1778
rect 3256 1678 3368 1738
rect 3256 1638 3292 1678
rect 3332 1638 3368 1678
rect 3256 1578 3368 1638
rect 3256 1538 3292 1578
rect 3332 1538 3368 1578
rect 3256 1478 3368 1538
rect 3256 1438 3292 1478
rect 3332 1438 3368 1478
rect 3256 1368 3368 1438
rect 3398 1778 3512 1848
rect 3398 1738 3436 1778
rect 3476 1738 3512 1778
rect 3398 1678 3512 1738
rect 3398 1638 3436 1678
rect 3476 1638 3512 1678
rect 3398 1578 3512 1638
rect 3398 1538 3436 1578
rect 3476 1538 3512 1578
rect 3398 1478 3512 1538
rect 3398 1438 3436 1478
rect 3476 1438 3512 1478
rect 3398 1368 3512 1438
rect 3542 1778 3656 1848
rect 3542 1738 3580 1778
rect 3620 1738 3656 1778
rect 3542 1678 3656 1738
rect 3542 1638 3580 1678
rect 3620 1638 3656 1678
rect 3542 1578 3656 1638
rect 3542 1538 3580 1578
rect 3620 1538 3656 1578
rect 3542 1478 3656 1538
rect 3542 1438 3580 1478
rect 3620 1438 3656 1478
rect 3542 1368 3656 1438
rect 3832 1778 3944 1848
rect 3832 1738 3868 1778
rect 3908 1738 3944 1778
rect 3832 1678 3944 1738
rect 3832 1638 3868 1678
rect 3908 1638 3944 1678
rect 3832 1578 3944 1638
rect 3832 1538 3868 1578
rect 3908 1538 3944 1578
rect 3832 1478 3944 1538
rect 3832 1438 3868 1478
rect 3908 1438 3944 1478
rect 3832 1368 3944 1438
rect 3974 1778 4088 1848
rect 3974 1738 4012 1778
rect 4052 1738 4088 1778
rect 3974 1678 4088 1738
rect 3974 1638 4012 1678
rect 4052 1638 4088 1678
rect 3974 1578 4088 1638
rect 3974 1538 4012 1578
rect 4052 1538 4088 1578
rect 3974 1478 4088 1538
rect 3974 1438 4012 1478
rect 4052 1438 4088 1478
rect 3974 1368 4088 1438
rect 4118 1778 4232 1848
rect 4118 1738 4156 1778
rect 4196 1738 4232 1778
rect 4118 1678 4232 1738
rect 4118 1638 4156 1678
rect 4196 1638 4232 1678
rect 4118 1578 4232 1638
rect 4118 1538 4156 1578
rect 4196 1538 4232 1578
rect 4118 1478 4232 1538
rect 4118 1438 4156 1478
rect 4196 1438 4232 1478
rect 4118 1368 4232 1438
rect 4408 1778 4520 1848
rect 4408 1738 4444 1778
rect 4484 1738 4520 1778
rect 4408 1678 4520 1738
rect 4408 1638 4444 1678
rect 4484 1638 4520 1678
rect 4408 1578 4520 1638
rect 4408 1538 4444 1578
rect 4484 1538 4520 1578
rect 4408 1478 4520 1538
rect 4408 1438 4444 1478
rect 4484 1438 4520 1478
rect 4408 1368 4520 1438
rect 4550 1778 4664 1848
rect 4550 1738 4588 1778
rect 4628 1738 4664 1778
rect 4550 1678 4664 1738
rect 4550 1638 4588 1678
rect 4628 1638 4664 1678
rect 4550 1578 4664 1638
rect 4550 1538 4588 1578
rect 4628 1538 4664 1578
rect 4550 1478 4664 1538
rect 4550 1438 4588 1478
rect 4628 1438 4664 1478
rect 4550 1368 4664 1438
rect 4694 1778 4808 1848
rect 4694 1738 4732 1778
rect 4772 1738 4808 1778
rect 4694 1678 4808 1738
rect 4694 1638 4732 1678
rect 4772 1638 4808 1678
rect 4694 1578 4808 1638
rect 4694 1538 4732 1578
rect 4772 1538 4808 1578
rect 4694 1478 4808 1538
rect 4694 1438 4732 1478
rect 4772 1438 4808 1478
rect 4694 1368 4808 1438
rect 4984 1778 5096 1848
rect 4984 1738 5020 1778
rect 5060 1738 5096 1778
rect 4984 1678 5096 1738
rect 4984 1638 5020 1678
rect 5060 1638 5096 1678
rect 4984 1578 5096 1638
rect 4984 1538 5020 1578
rect 5060 1538 5096 1578
rect 4984 1478 5096 1538
rect 4984 1438 5020 1478
rect 5060 1438 5096 1478
rect 4984 1368 5096 1438
rect 5126 1778 5240 1848
rect 5126 1738 5164 1778
rect 5204 1738 5240 1778
rect 5126 1678 5240 1738
rect 5126 1638 5164 1678
rect 5204 1638 5240 1678
rect 5126 1578 5240 1638
rect 5126 1538 5164 1578
rect 5204 1538 5240 1578
rect 5126 1478 5240 1538
rect 5126 1438 5164 1478
rect 5204 1438 5240 1478
rect 5126 1368 5240 1438
rect 5270 1778 5384 1848
rect 5270 1738 5308 1778
rect 5348 1738 5384 1778
rect 5270 1678 5384 1738
rect 5270 1638 5308 1678
rect 5348 1638 5384 1678
rect 5270 1578 5384 1638
rect 5270 1538 5308 1578
rect 5348 1538 5384 1578
rect 5270 1478 5384 1538
rect 5270 1438 5308 1478
rect 5348 1438 5384 1478
rect 5270 1368 5384 1438
rect 5848 1778 5960 1848
rect 5848 1738 5884 1778
rect 5924 1738 5960 1778
rect 5848 1678 5960 1738
rect 5848 1638 5884 1678
rect 5924 1638 5960 1678
rect 5848 1578 5960 1638
rect 5848 1538 5884 1578
rect 5924 1538 5960 1578
rect 5848 1478 5960 1538
rect 5848 1438 5884 1478
rect 5924 1438 5960 1478
rect 5848 1368 5960 1438
rect 5990 1778 6104 1848
rect 5990 1738 6028 1778
rect 6068 1738 6104 1778
rect 5990 1678 6104 1738
rect 5990 1638 6028 1678
rect 6068 1638 6104 1678
rect 5990 1578 6104 1638
rect 5990 1538 6028 1578
rect 6068 1538 6104 1578
rect 5990 1478 6104 1538
rect 5990 1438 6028 1478
rect 6068 1438 6104 1478
rect 5990 1368 6104 1438
rect 6134 1778 6248 1848
rect 6134 1738 6172 1778
rect 6212 1738 6248 1778
rect 6134 1678 6248 1738
rect 6134 1638 6172 1678
rect 6212 1638 6248 1678
rect 6134 1578 6248 1638
rect 6134 1538 6172 1578
rect 6212 1538 6248 1578
rect 6134 1478 6248 1538
rect 6134 1438 6172 1478
rect 6212 1438 6248 1478
rect 6134 1368 6248 1438
<< ndiffc >>
rect 124 558 164 598
rect 124 458 164 498
rect 268 558 308 598
rect 268 458 308 498
rect 412 558 452 598
rect 412 458 452 498
rect 700 558 740 598
rect 700 458 740 498
rect 844 558 884 598
rect 844 458 884 498
rect 988 558 1028 598
rect 988 458 1028 498
rect 1276 558 1316 598
rect 1276 458 1316 498
rect 1420 558 1460 598
rect 1420 458 1460 498
rect 1564 558 1604 598
rect 1564 458 1604 498
rect 1852 558 1892 598
rect 1852 458 1892 498
rect 1996 558 2036 598
rect 1996 458 2036 498
rect 2140 558 2180 598
rect 2140 458 2180 498
rect 2428 558 2468 598
rect 2428 458 2468 498
rect 2572 558 2612 598
rect 2572 458 2612 498
rect 2716 558 2756 598
rect 2716 458 2756 498
rect 3292 558 3332 598
rect 3292 458 3332 498
rect 3436 558 3476 598
rect 3436 458 3476 498
rect 3580 558 3620 598
rect 3580 458 3620 498
rect 3868 558 3908 598
rect 3868 458 3908 498
rect 4012 558 4052 598
rect 4012 458 4052 498
rect 4156 558 4196 598
rect 4156 458 4196 498
rect 4444 558 4484 598
rect 4444 458 4484 498
rect 4588 558 4628 598
rect 4588 458 4628 498
rect 4732 558 4772 598
rect 4732 458 4772 498
rect 5020 558 5060 598
rect 5020 458 5060 498
rect 5164 558 5204 598
rect 5164 458 5204 498
rect 5308 558 5348 598
rect 5308 458 5348 498
rect 5884 558 5924 598
rect 5884 458 5924 498
rect 6028 558 6068 598
rect 6028 458 6068 498
rect 6172 558 6212 598
rect 6172 458 6212 498
<< pdiffc >>
rect 124 1738 164 1778
rect 124 1638 164 1678
rect 124 1538 164 1578
rect 124 1438 164 1478
rect 268 1738 308 1778
rect 268 1638 308 1678
rect 268 1538 308 1578
rect 268 1438 308 1478
rect 412 1738 452 1778
rect 412 1638 452 1678
rect 412 1538 452 1578
rect 412 1438 452 1478
rect 700 1738 740 1778
rect 700 1638 740 1678
rect 700 1538 740 1578
rect 700 1438 740 1478
rect 844 1738 884 1778
rect 844 1638 884 1678
rect 844 1538 884 1578
rect 844 1438 884 1478
rect 988 1738 1028 1778
rect 988 1638 1028 1678
rect 988 1538 1028 1578
rect 988 1438 1028 1478
rect 1276 1738 1316 1778
rect 1276 1638 1316 1678
rect 1276 1538 1316 1578
rect 1276 1438 1316 1478
rect 1420 1738 1460 1778
rect 1420 1638 1460 1678
rect 1420 1538 1460 1578
rect 1420 1438 1460 1478
rect 1564 1738 1604 1778
rect 1564 1638 1604 1678
rect 1564 1538 1604 1578
rect 1564 1438 1604 1478
rect 1852 1738 1892 1778
rect 1852 1638 1892 1678
rect 1852 1538 1892 1578
rect 1852 1438 1892 1478
rect 1996 1738 2036 1778
rect 1996 1638 2036 1678
rect 1996 1538 2036 1578
rect 1996 1438 2036 1478
rect 2140 1738 2180 1778
rect 2140 1638 2180 1678
rect 2140 1538 2180 1578
rect 2140 1438 2180 1478
rect 2428 1738 2468 1778
rect 2428 1638 2468 1678
rect 2428 1538 2468 1578
rect 2428 1438 2468 1478
rect 2572 1738 2612 1778
rect 2572 1638 2612 1678
rect 2572 1538 2612 1578
rect 2572 1438 2612 1478
rect 2716 1738 2756 1778
rect 2716 1638 2756 1678
rect 2716 1538 2756 1578
rect 2716 1438 2756 1478
rect 3292 1738 3332 1778
rect 3292 1638 3332 1678
rect 3292 1538 3332 1578
rect 3292 1438 3332 1478
rect 3436 1738 3476 1778
rect 3436 1638 3476 1678
rect 3436 1538 3476 1578
rect 3436 1438 3476 1478
rect 3580 1738 3620 1778
rect 3580 1638 3620 1678
rect 3580 1538 3620 1578
rect 3580 1438 3620 1478
rect 3868 1738 3908 1778
rect 3868 1638 3908 1678
rect 3868 1538 3908 1578
rect 3868 1438 3908 1478
rect 4012 1738 4052 1778
rect 4012 1638 4052 1678
rect 4012 1538 4052 1578
rect 4012 1438 4052 1478
rect 4156 1738 4196 1778
rect 4156 1638 4196 1678
rect 4156 1538 4196 1578
rect 4156 1438 4196 1478
rect 4444 1738 4484 1778
rect 4444 1638 4484 1678
rect 4444 1538 4484 1578
rect 4444 1438 4484 1478
rect 4588 1738 4628 1778
rect 4588 1638 4628 1678
rect 4588 1538 4628 1578
rect 4588 1438 4628 1478
rect 4732 1738 4772 1778
rect 4732 1638 4772 1678
rect 4732 1538 4772 1578
rect 4732 1438 4772 1478
rect 5020 1738 5060 1778
rect 5020 1638 5060 1678
rect 5020 1538 5060 1578
rect 5020 1438 5060 1478
rect 5164 1738 5204 1778
rect 5164 1638 5204 1678
rect 5164 1538 5204 1578
rect 5164 1438 5204 1478
rect 5308 1738 5348 1778
rect 5308 1638 5348 1678
rect 5308 1538 5348 1578
rect 5308 1438 5348 1478
rect 5884 1738 5924 1778
rect 5884 1638 5924 1678
rect 5884 1538 5924 1578
rect 5884 1438 5924 1478
rect 6028 1738 6068 1778
rect 6028 1638 6068 1678
rect 6028 1538 6068 1578
rect 6028 1438 6068 1478
rect 6172 1738 6212 1778
rect 6172 1638 6212 1678
rect 6172 1538 6212 1578
rect 6172 1438 6212 1478
<< psubdiff >>
rect 5552 592 5760 642
rect 5552 450 5600 592
rect 5710 450 5760 592
rect 5552 406 5760 450
<< nsubdiff >>
rect 5472 1694 5760 1796
rect 5472 1450 5556 1694
rect 5682 1450 5760 1694
rect 5472 1390 5760 1450
<< psubdiffcont >>
rect 5600 450 5710 592
<< nsubdiffcont >>
rect 5556 1450 5682 1694
<< poly >>
rect 200 1848 230 1884
rect 344 1848 374 1884
rect 776 1848 806 1884
rect 920 1848 950 1884
rect 1352 1848 1382 1884
rect 1496 1848 1526 1884
rect 1928 1848 1958 1884
rect 2072 1848 2102 1884
rect 2504 1848 2534 1884
rect 2648 1848 2678 1884
rect 3368 1848 3398 1884
rect 3512 1848 3542 1884
rect 3944 1848 3974 1884
rect 4088 1848 4118 1884
rect 4520 1848 4550 1884
rect 4664 1848 4694 1884
rect 5096 1848 5126 1884
rect 5240 1848 5270 1884
rect 5960 1848 5990 1884
rect 6104 1848 6134 1884
rect 200 1332 230 1368
rect 344 1332 374 1368
rect 200 1313 374 1332
rect 200 1279 220 1313
rect 254 1279 328 1313
rect 362 1279 374 1313
rect 200 1260 374 1279
rect 776 1332 806 1368
rect 920 1332 950 1368
rect 776 1313 950 1332
rect 776 1279 796 1313
rect 830 1279 904 1313
rect 938 1279 950 1313
rect 776 1260 950 1279
rect 1352 1332 1382 1368
rect 1496 1332 1526 1368
rect 1352 1313 1526 1332
rect 1352 1279 1372 1313
rect 1406 1279 1480 1313
rect 1514 1279 1526 1313
rect 1352 1260 1526 1279
rect 1928 1332 1958 1368
rect 2072 1332 2102 1368
rect 2504 1332 2534 1368
rect 1928 1313 2102 1332
rect 1928 1279 1948 1313
rect 1982 1279 2056 1313
rect 2090 1279 2102 1313
rect 1928 1260 2102 1279
rect 2414 1314 2534 1332
rect 2414 1278 2436 1314
rect 2472 1278 2534 1314
rect 2414 1260 2534 1278
rect 2648 1332 2678 1368
rect 3368 1332 3398 1368
rect 3512 1332 3542 1368
rect 2648 1314 2768 1332
rect 2648 1278 2720 1314
rect 2756 1278 2768 1314
rect 2648 1260 2768 1278
rect 3368 1313 3542 1332
rect 3368 1279 3388 1313
rect 3422 1279 3496 1313
rect 3530 1279 3542 1313
rect 3368 1260 3542 1279
rect 3944 1332 3974 1368
rect 4088 1332 4118 1368
rect 3944 1313 4118 1332
rect 3944 1279 3964 1313
rect 3998 1279 4072 1313
rect 4106 1279 4118 1313
rect 3944 1260 4118 1279
rect 4520 1332 4550 1368
rect 4664 1332 4694 1368
rect 5096 1332 5126 1368
rect 4520 1313 4694 1332
rect 4520 1279 4540 1313
rect 4574 1279 4648 1313
rect 4682 1279 4694 1313
rect 4520 1260 4694 1279
rect 5006 1314 5126 1332
rect 5006 1278 5028 1314
rect 5064 1278 5126 1314
rect 5006 1260 5126 1278
rect 5240 1332 5270 1368
rect 5960 1332 5990 1368
rect 6104 1332 6134 1368
rect 5240 1314 5360 1332
rect 5240 1278 5312 1314
rect 5348 1278 5360 1314
rect 5240 1260 5360 1278
rect 5960 1313 6134 1332
rect 5960 1279 5980 1313
rect 6014 1279 6088 1313
rect 6122 1279 6134 1313
rect 5960 1260 6134 1279
rect 200 737 374 756
rect 200 703 220 737
rect 254 703 328 737
rect 362 703 374 737
rect 200 684 374 703
rect 200 648 230 684
rect 344 648 374 684
rect 776 737 950 756
rect 776 703 796 737
rect 830 703 904 737
rect 938 703 950 737
rect 776 684 950 703
rect 776 648 806 684
rect 920 648 950 684
rect 1352 737 1526 756
rect 1352 703 1372 737
rect 1406 703 1480 737
rect 1514 703 1526 737
rect 1352 684 1526 703
rect 1352 648 1382 684
rect 1496 648 1526 684
rect 1928 737 2102 756
rect 1928 703 1948 737
rect 1982 703 2056 737
rect 2090 703 2102 737
rect 1928 684 2102 703
rect 2414 738 2534 756
rect 2414 702 2436 738
rect 2472 702 2534 738
rect 2414 684 2534 702
rect 1928 648 1958 684
rect 2072 648 2102 684
rect 2504 648 2534 684
rect 2648 738 2768 756
rect 2648 702 2714 738
rect 2750 702 2768 738
rect 2648 684 2768 702
rect 3368 737 3542 756
rect 3368 703 3388 737
rect 3422 703 3496 737
rect 3530 703 3542 737
rect 3368 684 3542 703
rect 2648 648 2678 684
rect 3368 648 3398 684
rect 3512 648 3542 684
rect 3944 737 4118 756
rect 3944 703 3964 737
rect 3998 703 4072 737
rect 4106 703 4118 737
rect 3944 684 4118 703
rect 3944 648 3974 684
rect 4088 648 4118 684
rect 4520 737 4694 756
rect 4520 703 4540 737
rect 4574 703 4648 737
rect 4682 703 4694 737
rect 4520 684 4694 703
rect 5006 738 5126 756
rect 5006 702 5028 738
rect 5064 702 5126 738
rect 5006 684 5126 702
rect 4520 648 4550 684
rect 4664 648 4694 684
rect 5096 648 5126 684
rect 5240 738 5360 756
rect 5240 702 5306 738
rect 5342 702 5360 738
rect 5240 684 5360 702
rect 5960 737 6134 756
rect 5960 703 5980 737
rect 6014 703 6088 737
rect 6122 703 6134 737
rect 5960 684 6134 703
rect 5240 648 5270 684
rect 5960 648 5990 684
rect 6104 648 6134 684
rect 200 372 230 408
rect 344 372 374 408
rect 776 372 806 408
rect 920 372 950 408
rect 1352 372 1382 408
rect 1496 372 1526 408
rect 1928 372 1958 408
rect 2072 372 2102 408
rect 2504 372 2534 408
rect 2648 372 2678 408
rect 3368 372 3398 408
rect 3512 372 3542 408
rect 3944 372 3974 408
rect 4088 372 4118 408
rect 4520 372 4550 408
rect 4664 372 4694 408
rect 5096 372 5126 408
rect 5240 372 5270 408
rect 5960 372 5990 408
rect 6104 372 6134 408
<< polycont >>
rect 220 1279 254 1313
rect 328 1279 362 1313
rect 796 1279 830 1313
rect 904 1279 938 1313
rect 1372 1279 1406 1313
rect 1480 1279 1514 1313
rect 1948 1279 1982 1313
rect 2056 1279 2090 1313
rect 2436 1278 2472 1314
rect 2720 1278 2756 1314
rect 3388 1279 3422 1313
rect 3496 1279 3530 1313
rect 3964 1279 3998 1313
rect 4072 1279 4106 1313
rect 4540 1279 4574 1313
rect 4648 1279 4682 1313
rect 5028 1278 5064 1314
rect 5312 1278 5348 1314
rect 5980 1279 6014 1313
rect 6088 1279 6122 1313
rect 220 703 254 737
rect 328 703 362 737
rect 796 703 830 737
rect 904 703 938 737
rect 1372 703 1406 737
rect 1480 703 1514 737
rect 1948 703 1982 737
rect 2056 703 2090 737
rect 2436 702 2472 738
rect 2714 702 2750 738
rect 3388 703 3422 737
rect 3496 703 3530 737
rect 3964 703 3998 737
rect 4072 703 4106 737
rect 4540 703 4574 737
rect 4648 703 4682 737
rect 5028 702 5064 738
rect 5306 702 5342 738
rect 5980 703 6014 737
rect 6088 703 6122 737
<< locali >>
rect 114 1778 174 1794
rect 114 1738 124 1778
rect 164 1738 174 1778
rect 114 1678 174 1738
rect 114 1638 124 1678
rect 164 1638 174 1678
rect 114 1578 174 1638
rect 114 1538 124 1578
rect 164 1538 174 1578
rect 114 1478 174 1538
rect 114 1438 124 1478
rect 164 1438 174 1478
rect 114 1422 174 1438
rect 258 1778 318 1794
rect 258 1738 268 1778
rect 308 1738 318 1778
rect 258 1678 318 1738
rect 258 1638 268 1678
rect 308 1638 318 1678
rect 258 1578 318 1638
rect 258 1538 268 1578
rect 308 1538 318 1578
rect 258 1478 318 1538
rect 258 1438 268 1478
rect 308 1438 318 1478
rect 258 1422 318 1438
rect 402 1778 462 1794
rect 402 1738 412 1778
rect 452 1738 462 1778
rect 402 1678 462 1738
rect 402 1638 412 1678
rect 452 1638 462 1678
rect 402 1578 462 1638
rect 402 1538 412 1578
rect 452 1538 462 1578
rect 402 1478 462 1538
rect 402 1438 412 1478
rect 452 1438 462 1478
rect 402 1422 462 1438
rect 690 1778 750 1794
rect 690 1738 700 1778
rect 740 1738 750 1778
rect 690 1678 750 1738
rect 690 1638 700 1678
rect 740 1638 750 1678
rect 690 1578 750 1638
rect 690 1538 700 1578
rect 740 1538 750 1578
rect 690 1478 750 1538
rect 690 1438 700 1478
rect 740 1438 750 1478
rect 690 1422 750 1438
rect 834 1778 894 1794
rect 834 1738 844 1778
rect 884 1738 894 1778
rect 834 1678 894 1738
rect 834 1638 844 1678
rect 884 1638 894 1678
rect 834 1578 894 1638
rect 834 1538 844 1578
rect 884 1538 894 1578
rect 834 1478 894 1538
rect 834 1438 844 1478
rect 884 1438 894 1478
rect 834 1422 894 1438
rect 978 1778 1038 1794
rect 978 1738 988 1778
rect 1028 1738 1038 1778
rect 978 1678 1038 1738
rect 978 1638 988 1678
rect 1028 1638 1038 1678
rect 978 1578 1038 1638
rect 978 1538 988 1578
rect 1028 1538 1038 1578
rect 978 1478 1038 1538
rect 978 1438 988 1478
rect 1028 1438 1038 1478
rect 978 1422 1038 1438
rect 1266 1778 1326 1794
rect 1266 1738 1276 1778
rect 1316 1738 1326 1778
rect 1266 1678 1326 1738
rect 1266 1638 1276 1678
rect 1316 1638 1326 1678
rect 1266 1578 1326 1638
rect 1266 1538 1276 1578
rect 1316 1538 1326 1578
rect 1266 1478 1326 1538
rect 1266 1438 1276 1478
rect 1316 1438 1326 1478
rect 1266 1422 1326 1438
rect 1410 1778 1470 1794
rect 1410 1738 1420 1778
rect 1460 1738 1470 1778
rect 1410 1678 1470 1738
rect 1410 1638 1420 1678
rect 1460 1638 1470 1678
rect 1410 1578 1470 1638
rect 1410 1538 1420 1578
rect 1460 1538 1470 1578
rect 1410 1478 1470 1538
rect 1410 1438 1420 1478
rect 1460 1438 1470 1478
rect 1410 1422 1470 1438
rect 1554 1778 1614 1794
rect 1554 1738 1564 1778
rect 1604 1738 1614 1778
rect 1554 1678 1614 1738
rect 1554 1638 1564 1678
rect 1604 1638 1614 1678
rect 1554 1578 1614 1638
rect 1554 1538 1564 1578
rect 1604 1538 1614 1578
rect 1554 1478 1614 1538
rect 1554 1438 1564 1478
rect 1604 1438 1614 1478
rect 1554 1422 1614 1438
rect 1842 1778 1902 1794
rect 1842 1738 1852 1778
rect 1892 1738 1902 1778
rect 1842 1678 1902 1738
rect 1842 1638 1852 1678
rect 1892 1638 1902 1678
rect 1842 1578 1902 1638
rect 1842 1538 1852 1578
rect 1892 1538 1902 1578
rect 1842 1478 1902 1538
rect 1842 1438 1852 1478
rect 1892 1438 1902 1478
rect 1842 1422 1902 1438
rect 1986 1778 2046 1794
rect 1986 1738 1996 1778
rect 2036 1738 2046 1778
rect 1986 1678 2046 1738
rect 1986 1638 1996 1678
rect 2036 1638 2046 1678
rect 1986 1578 2046 1638
rect 1986 1538 1996 1578
rect 2036 1538 2046 1578
rect 1986 1478 2046 1538
rect 1986 1438 1996 1478
rect 2036 1438 2046 1478
rect 1986 1422 2046 1438
rect 2130 1778 2190 1794
rect 2130 1738 2140 1778
rect 2180 1738 2190 1778
rect 2130 1678 2190 1738
rect 2130 1638 2140 1678
rect 2180 1638 2190 1678
rect 2130 1578 2190 1638
rect 2130 1538 2140 1578
rect 2180 1538 2190 1578
rect 2130 1478 2190 1538
rect 2130 1438 2140 1478
rect 2180 1438 2190 1478
rect 2130 1422 2190 1438
rect 2418 1778 2478 1794
rect 2418 1738 2428 1778
rect 2468 1738 2478 1778
rect 2418 1678 2478 1738
rect 2418 1638 2428 1678
rect 2468 1638 2478 1678
rect 2418 1578 2478 1638
rect 2418 1538 2428 1578
rect 2468 1538 2478 1578
rect 2418 1478 2478 1538
rect 2418 1438 2428 1478
rect 2468 1438 2478 1478
rect 2418 1422 2478 1438
rect 2562 1778 2622 1794
rect 2562 1738 2572 1778
rect 2612 1738 2622 1778
rect 2562 1678 2622 1738
rect 2562 1638 2572 1678
rect 2612 1638 2622 1678
rect 2562 1578 2622 1638
rect 2562 1538 2572 1578
rect 2612 1538 2622 1578
rect 2562 1478 2622 1538
rect 2562 1438 2572 1478
rect 2612 1438 2622 1478
rect 2562 1422 2622 1438
rect 2706 1778 2766 1794
rect 2706 1738 2716 1778
rect 2756 1738 2766 1778
rect 2706 1678 2766 1738
rect 2706 1638 2716 1678
rect 2756 1638 2766 1678
rect 2706 1578 2766 1638
rect 2706 1538 2716 1578
rect 2756 1538 2766 1578
rect 2706 1478 2766 1538
rect 2706 1438 2716 1478
rect 2756 1438 2766 1478
rect 2706 1422 2766 1438
rect 3282 1778 3342 1794
rect 3282 1738 3292 1778
rect 3332 1738 3342 1778
rect 3282 1678 3342 1738
rect 3282 1638 3292 1678
rect 3332 1638 3342 1678
rect 3282 1578 3342 1638
rect 3282 1538 3292 1578
rect 3332 1538 3342 1578
rect 3282 1478 3342 1538
rect 3282 1438 3292 1478
rect 3332 1438 3342 1478
rect 3282 1422 3342 1438
rect 3426 1778 3486 1794
rect 3426 1738 3436 1778
rect 3476 1738 3486 1778
rect 3426 1678 3486 1738
rect 3426 1638 3436 1678
rect 3476 1638 3486 1678
rect 3426 1578 3486 1638
rect 3426 1538 3436 1578
rect 3476 1538 3486 1578
rect 3426 1478 3486 1538
rect 3426 1438 3436 1478
rect 3476 1438 3486 1478
rect 3426 1422 3486 1438
rect 3570 1778 3630 1794
rect 3570 1738 3580 1778
rect 3620 1738 3630 1778
rect 3570 1678 3630 1738
rect 3570 1638 3580 1678
rect 3620 1638 3630 1678
rect 3570 1578 3630 1638
rect 3570 1538 3580 1578
rect 3620 1538 3630 1578
rect 3570 1478 3630 1538
rect 3570 1438 3580 1478
rect 3620 1438 3630 1478
rect 3570 1422 3630 1438
rect 3858 1778 3918 1794
rect 3858 1738 3868 1778
rect 3908 1738 3918 1778
rect 3858 1678 3918 1738
rect 3858 1638 3868 1678
rect 3908 1638 3918 1678
rect 3858 1578 3918 1638
rect 3858 1538 3868 1578
rect 3908 1538 3918 1578
rect 3858 1478 3918 1538
rect 3858 1438 3868 1478
rect 3908 1438 3918 1478
rect 3858 1422 3918 1438
rect 4002 1778 4062 1794
rect 4002 1738 4012 1778
rect 4052 1738 4062 1778
rect 4002 1678 4062 1738
rect 4002 1638 4012 1678
rect 4052 1638 4062 1678
rect 4002 1578 4062 1638
rect 4002 1538 4012 1578
rect 4052 1538 4062 1578
rect 4002 1478 4062 1538
rect 4002 1438 4012 1478
rect 4052 1438 4062 1478
rect 4002 1422 4062 1438
rect 4146 1778 4206 1794
rect 4146 1738 4156 1778
rect 4196 1738 4206 1778
rect 4146 1678 4206 1738
rect 4146 1638 4156 1678
rect 4196 1638 4206 1678
rect 4146 1578 4206 1638
rect 4146 1538 4156 1578
rect 4196 1538 4206 1578
rect 4146 1478 4206 1538
rect 4146 1438 4156 1478
rect 4196 1438 4206 1478
rect 4146 1422 4206 1438
rect 4434 1778 4494 1794
rect 4434 1738 4444 1778
rect 4484 1738 4494 1778
rect 4434 1678 4494 1738
rect 4434 1638 4444 1678
rect 4484 1638 4494 1678
rect 4434 1578 4494 1638
rect 4434 1538 4444 1578
rect 4484 1538 4494 1578
rect 4434 1478 4494 1538
rect 4434 1438 4444 1478
rect 4484 1438 4494 1478
rect 4434 1422 4494 1438
rect 4578 1778 4638 1794
rect 4578 1738 4588 1778
rect 4628 1738 4638 1778
rect 4578 1678 4638 1738
rect 4578 1638 4588 1678
rect 4628 1638 4638 1678
rect 4578 1578 4638 1638
rect 4578 1538 4588 1578
rect 4628 1538 4638 1578
rect 4578 1478 4638 1538
rect 4578 1438 4588 1478
rect 4628 1438 4638 1478
rect 4578 1422 4638 1438
rect 4722 1778 4782 1794
rect 4722 1738 4732 1778
rect 4772 1738 4782 1778
rect 4722 1678 4782 1738
rect 4722 1638 4732 1678
rect 4772 1638 4782 1678
rect 4722 1578 4782 1638
rect 4722 1538 4732 1578
rect 4772 1538 4782 1578
rect 4722 1478 4782 1538
rect 4722 1438 4732 1478
rect 4772 1438 4782 1478
rect 4722 1422 4782 1438
rect 5010 1778 5070 1794
rect 5010 1738 5020 1778
rect 5060 1738 5070 1778
rect 5010 1678 5070 1738
rect 5010 1638 5020 1678
rect 5060 1638 5070 1678
rect 5010 1578 5070 1638
rect 5010 1538 5020 1578
rect 5060 1538 5070 1578
rect 5010 1478 5070 1538
rect 5010 1438 5020 1478
rect 5060 1438 5070 1478
rect 5010 1422 5070 1438
rect 5154 1778 5214 1794
rect 5154 1738 5164 1778
rect 5204 1738 5214 1778
rect 5154 1678 5214 1738
rect 5154 1638 5164 1678
rect 5204 1638 5214 1678
rect 5154 1578 5214 1638
rect 5154 1538 5164 1578
rect 5204 1538 5214 1578
rect 5154 1478 5214 1538
rect 5154 1438 5164 1478
rect 5204 1438 5214 1478
rect 5154 1422 5214 1438
rect 5298 1778 5358 1794
rect 5298 1738 5308 1778
rect 5348 1738 5358 1778
rect 5298 1678 5358 1738
rect 5298 1638 5308 1678
rect 5348 1638 5358 1678
rect 5298 1578 5358 1638
rect 5298 1538 5308 1578
rect 5348 1538 5358 1578
rect 5298 1478 5358 1538
rect 5298 1438 5308 1478
rect 5348 1438 5358 1478
rect 5298 1422 5358 1438
rect 5472 1694 5760 1796
rect 5472 1450 5556 1694
rect 5682 1450 5760 1694
rect 5472 1390 5760 1450
rect 5874 1778 5934 1794
rect 5874 1738 5884 1778
rect 5924 1738 5934 1778
rect 5874 1678 5934 1738
rect 5874 1638 5884 1678
rect 5924 1638 5934 1678
rect 5874 1578 5934 1638
rect 5874 1538 5884 1578
rect 5924 1538 5934 1578
rect 5874 1478 5934 1538
rect 5874 1438 5884 1478
rect 5924 1438 5934 1478
rect 5874 1422 5934 1438
rect 6018 1778 6078 1794
rect 6018 1738 6028 1778
rect 6068 1738 6078 1778
rect 6018 1678 6078 1738
rect 6018 1638 6028 1678
rect 6068 1638 6078 1678
rect 6018 1578 6078 1638
rect 6018 1538 6028 1578
rect 6068 1538 6078 1578
rect 6018 1478 6078 1538
rect 6018 1438 6028 1478
rect 6068 1438 6078 1478
rect 6018 1422 6078 1438
rect 6162 1778 6222 1794
rect 6162 1738 6172 1778
rect 6212 1738 6222 1778
rect 6162 1678 6222 1738
rect 6162 1638 6172 1678
rect 6212 1638 6222 1678
rect 6162 1578 6222 1638
rect 6162 1538 6172 1578
rect 6212 1538 6222 1578
rect 6162 1478 6222 1538
rect 6162 1438 6172 1478
rect 6212 1438 6222 1478
rect 6162 1422 6222 1438
rect 200 1313 374 1332
rect 200 1279 220 1313
rect 254 1279 328 1313
rect 362 1279 374 1313
rect 200 1260 374 1279
rect 776 1313 950 1332
rect 776 1279 796 1313
rect 830 1279 904 1313
rect 938 1279 950 1313
rect 776 1260 950 1279
rect 1352 1313 1526 1332
rect 1352 1279 1372 1313
rect 1406 1279 1480 1313
rect 1514 1279 1526 1313
rect 1352 1260 1526 1279
rect 1928 1313 2102 1332
rect 1928 1279 1948 1313
rect 1982 1279 2056 1313
rect 2090 1279 2102 1313
rect 1928 1260 2102 1279
rect 2414 1314 2504 1332
rect 2414 1278 2436 1314
rect 2472 1278 2504 1314
rect 2414 1260 2504 1278
rect 2678 1314 2768 1332
rect 2678 1278 2720 1314
rect 2756 1278 2768 1314
rect 2678 1260 2768 1278
rect 3368 1313 3542 1332
rect 3368 1279 3388 1313
rect 3422 1279 3496 1313
rect 3530 1279 3542 1313
rect 3368 1260 3542 1279
rect 3944 1313 4118 1332
rect 3944 1279 3964 1313
rect 3998 1279 4072 1313
rect 4106 1279 4118 1313
rect 3944 1260 4118 1279
rect 4520 1313 4694 1332
rect 4520 1279 4540 1313
rect 4574 1279 4648 1313
rect 4682 1279 4694 1313
rect 4520 1260 4694 1279
rect 5006 1314 5096 1332
rect 5006 1278 5028 1314
rect 5064 1278 5096 1314
rect 5006 1260 5096 1278
rect 5270 1314 5360 1332
rect 5270 1278 5312 1314
rect 5348 1278 5360 1314
rect 5270 1260 5360 1278
rect 5960 1313 6134 1332
rect 5960 1279 5980 1313
rect 6014 1279 6088 1313
rect 6122 1279 6134 1313
rect 5960 1260 6134 1279
rect 200 737 374 756
rect 200 703 220 737
rect 254 703 328 737
rect 362 703 374 737
rect 200 684 374 703
rect 776 737 950 756
rect 776 703 796 737
rect 830 703 904 737
rect 938 703 950 737
rect 776 684 950 703
rect 1352 737 1526 756
rect 1352 703 1372 737
rect 1406 703 1480 737
rect 1514 703 1526 737
rect 1352 684 1526 703
rect 1928 737 2102 756
rect 1928 703 1948 737
rect 1982 703 2056 737
rect 2090 703 2102 737
rect 1928 684 2102 703
rect 2414 738 2504 756
rect 2414 702 2436 738
rect 2472 702 2504 738
rect 2414 684 2504 702
rect 2678 738 2768 756
rect 2678 702 2714 738
rect 2750 702 2768 738
rect 2678 684 2768 702
rect 3368 737 3542 756
rect 3368 703 3388 737
rect 3422 703 3496 737
rect 3530 703 3542 737
rect 3368 684 3542 703
rect 3944 737 4118 756
rect 3944 703 3964 737
rect 3998 703 4072 737
rect 4106 703 4118 737
rect 3944 684 4118 703
rect 4520 737 4694 756
rect 4520 703 4540 737
rect 4574 703 4648 737
rect 4682 703 4694 737
rect 4520 684 4694 703
rect 5006 738 5096 756
rect 5006 702 5028 738
rect 5064 702 5096 738
rect 5006 684 5096 702
rect 5270 738 5360 756
rect 5270 702 5306 738
rect 5342 702 5360 738
rect 5270 684 5360 702
rect 5960 737 6134 756
rect 5960 703 5980 737
rect 6014 703 6088 737
rect 6122 703 6134 737
rect 5960 684 6134 703
rect 114 598 174 614
rect 114 558 124 598
rect 164 558 174 598
rect 114 498 174 558
rect 114 458 124 498
rect 164 458 174 498
rect 114 442 174 458
rect 258 598 318 614
rect 258 558 268 598
rect 308 558 318 598
rect 258 498 318 558
rect 258 458 268 498
rect 308 458 318 498
rect 258 442 318 458
rect 402 598 462 614
rect 402 558 412 598
rect 452 558 462 598
rect 402 498 462 558
rect 402 458 412 498
rect 452 458 462 498
rect 402 442 462 458
rect 690 598 750 614
rect 690 558 700 598
rect 740 558 750 598
rect 690 498 750 558
rect 690 458 700 498
rect 740 458 750 498
rect 690 442 750 458
rect 834 598 894 614
rect 834 558 844 598
rect 884 558 894 598
rect 834 498 894 558
rect 834 458 844 498
rect 884 458 894 498
rect 834 442 894 458
rect 978 598 1038 614
rect 978 558 988 598
rect 1028 558 1038 598
rect 978 498 1038 558
rect 978 458 988 498
rect 1028 458 1038 498
rect 978 442 1038 458
rect 1266 598 1326 614
rect 1266 558 1276 598
rect 1316 558 1326 598
rect 1266 498 1326 558
rect 1266 458 1276 498
rect 1316 458 1326 498
rect 1266 442 1326 458
rect 1410 598 1470 614
rect 1410 558 1420 598
rect 1460 558 1470 598
rect 1410 498 1470 558
rect 1410 458 1420 498
rect 1460 458 1470 498
rect 1410 442 1470 458
rect 1554 598 1614 614
rect 1554 558 1564 598
rect 1604 558 1614 598
rect 1554 498 1614 558
rect 1554 458 1564 498
rect 1604 458 1614 498
rect 1554 442 1614 458
rect 1842 598 1902 614
rect 1842 558 1852 598
rect 1892 558 1902 598
rect 1842 498 1902 558
rect 1842 458 1852 498
rect 1892 458 1902 498
rect 1842 442 1902 458
rect 1986 598 2046 614
rect 1986 558 1996 598
rect 2036 558 2046 598
rect 1986 498 2046 558
rect 1986 458 1996 498
rect 2036 458 2046 498
rect 1986 442 2046 458
rect 2130 598 2190 614
rect 2130 558 2140 598
rect 2180 558 2190 598
rect 2130 498 2190 558
rect 2130 458 2140 498
rect 2180 458 2190 498
rect 2130 442 2190 458
rect 2418 598 2478 614
rect 2418 558 2428 598
rect 2468 558 2478 598
rect 2418 498 2478 558
rect 2418 458 2428 498
rect 2468 458 2478 498
rect 2418 442 2478 458
rect 2562 598 2622 614
rect 2562 558 2572 598
rect 2612 558 2622 598
rect 2562 498 2622 558
rect 2562 458 2572 498
rect 2612 458 2622 498
rect 2562 442 2622 458
rect 2706 598 2766 614
rect 2706 558 2716 598
rect 2756 558 2766 598
rect 2706 498 2766 558
rect 2706 458 2716 498
rect 2756 458 2766 498
rect 2706 442 2766 458
rect 3282 598 3342 614
rect 3282 558 3292 598
rect 3332 558 3342 598
rect 3282 498 3342 558
rect 3282 458 3292 498
rect 3332 458 3342 498
rect 3282 442 3342 458
rect 3426 598 3486 614
rect 3426 558 3436 598
rect 3476 558 3486 598
rect 3426 498 3486 558
rect 3426 458 3436 498
rect 3476 458 3486 498
rect 3426 442 3486 458
rect 3570 598 3630 614
rect 3570 558 3580 598
rect 3620 558 3630 598
rect 3570 498 3630 558
rect 3570 458 3580 498
rect 3620 458 3630 498
rect 3570 442 3630 458
rect 3858 598 3918 614
rect 3858 558 3868 598
rect 3908 558 3918 598
rect 3858 498 3918 558
rect 3858 458 3868 498
rect 3908 458 3918 498
rect 3858 442 3918 458
rect 4002 598 4062 614
rect 4002 558 4012 598
rect 4052 558 4062 598
rect 4002 498 4062 558
rect 4002 458 4012 498
rect 4052 458 4062 498
rect 4002 442 4062 458
rect 4146 598 4206 614
rect 4146 558 4156 598
rect 4196 558 4206 598
rect 4146 498 4206 558
rect 4146 458 4156 498
rect 4196 458 4206 498
rect 4146 442 4206 458
rect 4434 598 4494 614
rect 4434 558 4444 598
rect 4484 558 4494 598
rect 4434 498 4494 558
rect 4434 458 4444 498
rect 4484 458 4494 498
rect 4434 442 4494 458
rect 4578 598 4638 614
rect 4578 558 4588 598
rect 4628 558 4638 598
rect 4578 498 4638 558
rect 4578 458 4588 498
rect 4628 458 4638 498
rect 4578 442 4638 458
rect 4722 598 4782 614
rect 4722 558 4732 598
rect 4772 558 4782 598
rect 4722 498 4782 558
rect 4722 458 4732 498
rect 4772 458 4782 498
rect 4722 442 4782 458
rect 5010 598 5070 614
rect 5010 558 5020 598
rect 5060 558 5070 598
rect 5010 498 5070 558
rect 5010 458 5020 498
rect 5060 458 5070 498
rect 5010 442 5070 458
rect 5154 598 5214 614
rect 5154 558 5164 598
rect 5204 558 5214 598
rect 5154 498 5214 558
rect 5154 458 5164 498
rect 5204 458 5214 498
rect 5154 442 5214 458
rect 5298 598 5358 614
rect 5298 558 5308 598
rect 5348 558 5358 598
rect 5298 498 5358 558
rect 5298 458 5308 498
rect 5348 458 5358 498
rect 5298 442 5358 458
rect 5552 592 5760 642
rect 5552 450 5600 592
rect 5710 450 5760 592
rect 5552 406 5760 450
rect 5874 598 5934 614
rect 5874 558 5884 598
rect 5924 558 5934 598
rect 5874 498 5934 558
rect 5874 458 5884 498
rect 5924 458 5934 498
rect 5874 442 5934 458
rect 6018 598 6078 614
rect 6018 558 6028 598
rect 6068 558 6078 598
rect 6018 498 6078 558
rect 6018 458 6028 498
rect 6068 458 6078 498
rect 6018 442 6078 458
rect 6162 598 6222 614
rect 6162 558 6172 598
rect 6212 558 6222 598
rect 6162 498 6222 558
rect 6162 458 6172 498
rect 6212 458 6222 498
rect 6162 442 6222 458
<< viali >>
rect 124 1738 164 1778
rect 124 1638 164 1678
rect 124 1538 164 1578
rect 124 1438 164 1478
rect 268 1738 308 1778
rect 268 1638 308 1678
rect 268 1538 308 1578
rect 268 1438 308 1478
rect 412 1738 452 1778
rect 412 1638 452 1678
rect 412 1538 452 1578
rect 412 1438 452 1478
rect 700 1738 740 1778
rect 700 1638 740 1678
rect 700 1538 740 1578
rect 700 1438 740 1478
rect 844 1738 884 1778
rect 844 1638 884 1678
rect 844 1538 884 1578
rect 844 1438 884 1478
rect 988 1738 1028 1778
rect 988 1638 1028 1678
rect 988 1538 1028 1578
rect 988 1438 1028 1478
rect 1276 1738 1316 1778
rect 1276 1638 1316 1678
rect 1276 1538 1316 1578
rect 1276 1438 1316 1478
rect 1420 1738 1460 1778
rect 1420 1638 1460 1678
rect 1420 1538 1460 1578
rect 1420 1438 1460 1478
rect 1564 1738 1604 1778
rect 1564 1638 1604 1678
rect 1564 1538 1604 1578
rect 1564 1438 1604 1478
rect 1852 1738 1892 1778
rect 1852 1638 1892 1678
rect 1852 1538 1892 1578
rect 1852 1438 1892 1478
rect 1996 1738 2036 1778
rect 1996 1638 2036 1678
rect 1996 1538 2036 1578
rect 1996 1438 2036 1478
rect 2140 1738 2180 1778
rect 2140 1638 2180 1678
rect 2140 1538 2180 1578
rect 2140 1438 2180 1478
rect 2428 1738 2468 1778
rect 2428 1638 2468 1678
rect 2428 1538 2468 1578
rect 2428 1438 2468 1478
rect 2572 1738 2612 1778
rect 2572 1638 2612 1678
rect 2572 1538 2612 1578
rect 2572 1438 2612 1478
rect 2716 1738 2756 1778
rect 2716 1638 2756 1678
rect 2716 1538 2756 1578
rect 2716 1438 2756 1478
rect 3292 1738 3332 1778
rect 3292 1638 3332 1678
rect 3292 1538 3332 1578
rect 3292 1438 3332 1478
rect 3436 1738 3476 1778
rect 3436 1638 3476 1678
rect 3436 1538 3476 1578
rect 3436 1438 3476 1478
rect 3580 1738 3620 1778
rect 3580 1638 3620 1678
rect 3580 1538 3620 1578
rect 3580 1438 3620 1478
rect 3868 1738 3908 1778
rect 3868 1638 3908 1678
rect 3868 1538 3908 1578
rect 3868 1438 3908 1478
rect 4012 1738 4052 1778
rect 4012 1638 4052 1678
rect 4012 1538 4052 1578
rect 4012 1438 4052 1478
rect 4156 1738 4196 1778
rect 4156 1638 4196 1678
rect 4156 1538 4196 1578
rect 4156 1438 4196 1478
rect 4444 1738 4484 1778
rect 4444 1638 4484 1678
rect 4444 1538 4484 1578
rect 4444 1438 4484 1478
rect 4588 1738 4628 1778
rect 4588 1638 4628 1678
rect 4588 1538 4628 1578
rect 4588 1438 4628 1478
rect 4732 1738 4772 1778
rect 4732 1638 4772 1678
rect 4732 1538 4772 1578
rect 4732 1438 4772 1478
rect 5020 1738 5060 1778
rect 5020 1638 5060 1678
rect 5020 1538 5060 1578
rect 5020 1438 5060 1478
rect 5164 1738 5204 1778
rect 5164 1638 5204 1678
rect 5164 1538 5204 1578
rect 5164 1438 5204 1478
rect 5308 1738 5348 1778
rect 5308 1638 5348 1678
rect 5308 1538 5348 1578
rect 5308 1438 5348 1478
rect 5572 1476 5652 1666
rect 5884 1738 5924 1778
rect 5884 1638 5924 1678
rect 5884 1538 5924 1578
rect 5884 1438 5924 1478
rect 6028 1738 6068 1778
rect 6028 1638 6068 1678
rect 6028 1538 6068 1578
rect 6028 1438 6068 1478
rect 6172 1738 6212 1778
rect 6172 1638 6212 1678
rect 6172 1538 6212 1578
rect 6172 1438 6212 1478
rect 220 1279 254 1313
rect 328 1279 362 1313
rect 796 1279 830 1313
rect 904 1279 938 1313
rect 1372 1279 1406 1313
rect 1480 1279 1514 1313
rect 1948 1279 1982 1313
rect 2056 1279 2090 1313
rect 2436 1278 2472 1314
rect 2720 1278 2756 1314
rect 3388 1279 3422 1313
rect 3496 1279 3530 1313
rect 3964 1279 3998 1313
rect 4072 1279 4106 1313
rect 4540 1279 4574 1313
rect 4648 1279 4682 1313
rect 5028 1278 5064 1314
rect 5312 1278 5348 1314
rect 5980 1279 6014 1313
rect 6088 1279 6122 1313
rect 220 703 254 737
rect 328 703 362 737
rect 796 703 830 737
rect 904 703 938 737
rect 1372 703 1406 737
rect 1480 703 1514 737
rect 1948 703 1982 737
rect 2056 703 2090 737
rect 2436 702 2472 738
rect 2714 702 2750 738
rect 3388 703 3422 737
rect 3496 703 3530 737
rect 3964 703 3998 737
rect 4072 703 4106 737
rect 4540 703 4574 737
rect 4648 703 4682 737
rect 5028 702 5064 738
rect 5306 702 5342 738
rect 5980 703 6014 737
rect 6088 703 6122 737
rect 124 558 164 598
rect 124 458 164 498
rect 268 558 308 598
rect 268 458 308 498
rect 412 558 452 598
rect 412 458 452 498
rect 700 558 740 598
rect 700 458 740 498
rect 844 558 884 598
rect 844 458 884 498
rect 988 558 1028 598
rect 988 458 1028 498
rect 1276 558 1316 598
rect 1276 458 1316 498
rect 1420 558 1460 598
rect 1420 458 1460 498
rect 1564 558 1604 598
rect 1564 458 1604 498
rect 1852 558 1892 598
rect 1852 458 1892 498
rect 1996 558 2036 598
rect 1996 458 2036 498
rect 2140 558 2180 598
rect 2140 458 2180 498
rect 2428 558 2468 598
rect 2428 458 2468 498
rect 2572 558 2612 598
rect 2572 458 2612 498
rect 2716 558 2756 598
rect 2716 458 2756 498
rect 3292 558 3332 598
rect 3292 458 3332 498
rect 3436 558 3476 598
rect 3436 458 3476 498
rect 3580 558 3620 598
rect 3580 458 3620 498
rect 3868 558 3908 598
rect 3868 458 3908 498
rect 4012 558 4052 598
rect 4012 458 4052 498
rect 4156 558 4196 598
rect 4156 458 4196 498
rect 4444 558 4484 598
rect 4444 458 4484 498
rect 4588 558 4628 598
rect 4588 458 4628 498
rect 4732 558 4772 598
rect 4732 458 4772 498
rect 5020 558 5060 598
rect 5020 458 5060 498
rect 5164 558 5204 598
rect 5164 458 5204 498
rect 5308 558 5348 598
rect 5308 458 5348 498
rect 5600 450 5710 592
rect 5884 558 5924 598
rect 5884 458 5924 498
rect 6028 558 6068 598
rect 6028 458 6068 498
rect 6172 558 6212 598
rect 6172 458 6212 498
<< metal1 >>
rect 114 2048 174 2056
rect 402 2048 462 2056
rect 690 2048 750 2056
rect 978 2048 1038 2056
rect 1266 2048 1326 2056
rect 1554 2048 1614 2056
rect 3282 2048 3342 2056
rect 3570 2048 3630 2056
rect 3858 2048 3918 2056
rect 4146 2048 4206 2056
rect 112 2042 176 2048
rect 112 1990 118 2042
rect 170 1990 176 2042
rect 112 1984 176 1990
rect 400 2042 464 2048
rect 400 1990 406 2042
rect 458 1990 464 2042
rect 400 1984 464 1990
rect 688 2042 752 2048
rect 688 1990 694 2042
rect 746 1990 752 2042
rect 688 1984 752 1990
rect 976 2042 1040 2048
rect 976 1990 982 2042
rect 1034 1990 1040 2042
rect 976 1984 1040 1990
rect 1264 2042 1328 2048
rect 1264 1990 1270 2042
rect 1322 1990 1328 2042
rect 1264 1984 1328 1990
rect 1552 2042 1616 2048
rect 1552 1990 1558 2042
rect 1610 1990 1616 2042
rect 1552 1984 1616 1990
rect 2416 2042 2480 2048
rect 2416 1990 2422 2042
rect 2474 1990 2480 2042
rect 2416 1984 2480 1990
rect 3280 2042 3344 2048
rect 3280 1990 3286 2042
rect 3338 1990 3344 2042
rect 3280 1984 3344 1990
rect 3568 2042 3632 2048
rect 3568 1990 3574 2042
rect 3626 1990 3632 2042
rect 3568 1984 3632 1990
rect 3856 2042 3920 2048
rect 3856 1990 3862 2042
rect 3914 1990 3920 2042
rect 3856 1984 3920 1990
rect 4144 2042 4208 2048
rect 4144 1990 4150 2042
rect 4202 1990 4208 2042
rect 4144 1984 4208 1990
rect 5008 2042 5072 2048
rect 5008 1990 5014 2042
rect 5066 1990 5072 2042
rect 5008 1984 5072 1990
rect 5538 2044 5708 2052
rect 5874 2048 5934 2056
rect 6162 2048 6222 2056
rect 114 1778 174 1984
rect 114 1738 124 1778
rect 164 1738 174 1778
rect 114 1678 174 1738
rect 114 1638 124 1678
rect 164 1638 174 1678
rect 114 1578 174 1638
rect 258 1778 318 1828
rect 258 1738 268 1778
rect 308 1738 318 1778
rect 258 1678 318 1738
rect 258 1638 268 1678
rect 308 1638 318 1678
rect 258 1616 318 1638
rect 402 1778 462 1984
rect 402 1738 412 1778
rect 452 1738 462 1778
rect 402 1678 462 1738
rect 402 1638 412 1678
rect 452 1638 462 1678
rect 114 1538 124 1578
rect 164 1538 174 1578
rect 256 1610 320 1616
rect 256 1558 262 1610
rect 314 1558 320 1610
rect 256 1552 268 1558
rect 114 1478 174 1538
rect 114 1438 124 1478
rect 164 1438 174 1478
rect 114 1422 174 1438
rect 258 1538 268 1552
rect 308 1552 320 1558
rect 402 1578 462 1638
rect 308 1538 318 1552
rect 258 1478 318 1538
rect 258 1438 268 1478
rect 308 1438 318 1478
rect 258 1422 318 1438
rect 402 1538 412 1578
rect 452 1538 462 1578
rect 402 1478 462 1538
rect 402 1438 412 1478
rect 452 1438 462 1478
rect 402 1422 462 1438
rect 690 1778 750 1984
rect 690 1738 700 1778
rect 740 1738 750 1778
rect 690 1678 750 1738
rect 690 1638 700 1678
rect 740 1638 750 1678
rect 690 1578 750 1638
rect 834 1778 894 1828
rect 834 1738 844 1778
rect 884 1738 894 1778
rect 834 1678 894 1738
rect 834 1638 844 1678
rect 884 1638 894 1678
rect 834 1616 894 1638
rect 978 1778 1038 1984
rect 978 1738 988 1778
rect 1028 1738 1038 1778
rect 978 1678 1038 1738
rect 978 1638 988 1678
rect 1028 1638 1038 1678
rect 690 1538 700 1578
rect 740 1538 750 1578
rect 832 1610 896 1616
rect 832 1558 838 1610
rect 890 1558 896 1610
rect 832 1552 844 1558
rect 690 1478 750 1538
rect 690 1438 700 1478
rect 740 1438 750 1478
rect 690 1422 750 1438
rect 834 1538 844 1552
rect 884 1552 896 1558
rect 978 1578 1038 1638
rect 884 1538 894 1552
rect 834 1478 894 1538
rect 834 1438 844 1478
rect 884 1438 894 1478
rect 834 1422 894 1438
rect 978 1538 988 1578
rect 1028 1538 1038 1578
rect 978 1478 1038 1538
rect 978 1438 988 1478
rect 1028 1438 1038 1478
rect 978 1422 1038 1438
rect 1266 1778 1326 1984
rect 1266 1738 1276 1778
rect 1316 1738 1326 1778
rect 1266 1678 1326 1738
rect 1266 1638 1276 1678
rect 1316 1638 1326 1678
rect 1266 1578 1326 1638
rect 1410 1778 1470 1828
rect 1410 1738 1420 1778
rect 1460 1738 1470 1778
rect 1410 1678 1470 1738
rect 1410 1638 1420 1678
rect 1460 1638 1470 1678
rect 1410 1616 1470 1638
rect 1554 1778 1614 1984
rect 1554 1738 1564 1778
rect 1604 1738 1614 1778
rect 1554 1678 1614 1738
rect 1554 1638 1564 1678
rect 1604 1638 1614 1678
rect 1266 1538 1276 1578
rect 1316 1538 1326 1578
rect 1408 1610 1472 1616
rect 1408 1558 1414 1610
rect 1466 1558 1472 1610
rect 1408 1552 1420 1558
rect 1266 1478 1326 1538
rect 1266 1438 1276 1478
rect 1316 1438 1326 1478
rect 1266 1422 1326 1438
rect 1410 1538 1420 1552
rect 1460 1552 1472 1558
rect 1554 1578 1614 1638
rect 1842 1778 1902 1828
rect 1842 1738 1852 1778
rect 1892 1738 1902 1778
rect 1986 1778 2046 1828
rect 1986 1760 1996 1778
rect 1842 1678 1902 1738
rect 1984 1754 1996 1760
rect 2036 1760 2046 1778
rect 2130 1778 2190 1828
rect 2036 1754 2048 1760
rect 1984 1702 1990 1754
rect 2042 1702 2048 1754
rect 1984 1696 2048 1702
rect 2130 1738 2140 1778
rect 2180 1738 2190 1778
rect 1842 1638 1852 1678
rect 1892 1638 1902 1678
rect 1842 1616 1902 1638
rect 1986 1678 2046 1696
rect 1986 1638 1996 1678
rect 2036 1638 2046 1678
rect 1460 1538 1470 1552
rect 1410 1478 1470 1538
rect 1410 1438 1420 1478
rect 1460 1438 1470 1478
rect 1410 1422 1470 1438
rect 1554 1538 1564 1578
rect 1604 1538 1614 1578
rect 1840 1610 1904 1616
rect 1840 1558 1846 1610
rect 1898 1558 1904 1610
rect 1840 1552 1852 1558
rect 1554 1478 1614 1538
rect 1554 1438 1564 1478
rect 1604 1438 1614 1478
rect 1554 1422 1614 1438
rect 1842 1538 1852 1552
rect 1892 1552 1904 1558
rect 1986 1578 2046 1638
rect 2130 1678 2190 1738
rect 2130 1638 2140 1678
rect 2180 1638 2190 1678
rect 2130 1616 2190 1638
rect 2418 1778 2478 1984
rect 2418 1738 2428 1778
rect 2468 1738 2478 1778
rect 2418 1678 2478 1738
rect 2418 1638 2428 1678
rect 2468 1638 2478 1678
rect 1892 1538 1902 1552
rect 1842 1478 1902 1538
rect 1842 1438 1852 1478
rect 1892 1438 1902 1478
rect 1842 1422 1902 1438
rect 1986 1538 1996 1578
rect 2036 1538 2046 1578
rect 2128 1610 2192 1616
rect 2128 1558 2134 1610
rect 2186 1558 2192 1610
rect 2128 1552 2140 1558
rect 1986 1478 2046 1538
rect 1986 1438 1996 1478
rect 2036 1438 2046 1478
rect 1986 1422 2046 1438
rect 2130 1538 2140 1552
rect 2180 1552 2192 1558
rect 2418 1578 2478 1638
rect 2180 1538 2190 1552
rect 2130 1478 2190 1538
rect 2130 1438 2140 1478
rect 2180 1438 2190 1478
rect 2130 1422 2190 1438
rect 2418 1538 2428 1578
rect 2468 1538 2478 1578
rect 2418 1478 2478 1538
rect 2418 1438 2428 1478
rect 2468 1438 2478 1478
rect 2418 1422 2478 1438
rect 2562 1778 2622 1828
rect 2562 1738 2572 1778
rect 2612 1738 2622 1778
rect 2706 1778 2766 1828
rect 2706 1760 2716 1778
rect 2562 1678 2622 1738
rect 2704 1754 2716 1760
rect 2756 1760 2766 1778
rect 3282 1778 3342 1984
rect 2756 1754 2768 1760
rect 2704 1702 2710 1754
rect 2762 1702 2768 1754
rect 2704 1696 2768 1702
rect 3282 1738 3292 1778
rect 3332 1738 3342 1778
rect 2562 1638 2572 1678
rect 2612 1638 2622 1678
rect 2562 1578 2622 1638
rect 2562 1538 2572 1578
rect 2612 1538 2622 1578
rect 2562 1478 2622 1538
rect 2562 1438 2572 1478
rect 2612 1438 2622 1478
rect 2562 1422 2622 1438
rect 2706 1678 2766 1696
rect 2706 1638 2716 1678
rect 2756 1638 2766 1678
rect 2706 1578 2766 1638
rect 2706 1538 2716 1578
rect 2756 1538 2766 1578
rect 2706 1478 2766 1538
rect 2706 1438 2716 1478
rect 2756 1438 2766 1478
rect 2706 1422 2766 1438
rect 3282 1678 3342 1738
rect 3282 1638 3292 1678
rect 3332 1638 3342 1678
rect 3282 1578 3342 1638
rect 3426 1778 3486 1828
rect 3426 1738 3436 1778
rect 3476 1738 3486 1778
rect 3426 1678 3486 1738
rect 3426 1638 3436 1678
rect 3476 1638 3486 1678
rect 3426 1616 3486 1638
rect 3570 1778 3630 1984
rect 3570 1738 3580 1778
rect 3620 1738 3630 1778
rect 3570 1678 3630 1738
rect 3570 1638 3580 1678
rect 3620 1638 3630 1678
rect 3282 1538 3292 1578
rect 3332 1538 3342 1578
rect 3424 1610 3488 1616
rect 3424 1558 3430 1610
rect 3482 1558 3488 1610
rect 3424 1552 3436 1558
rect 3282 1478 3342 1538
rect 3282 1438 3292 1478
rect 3332 1438 3342 1478
rect 3282 1422 3342 1438
rect 3426 1538 3436 1552
rect 3476 1552 3488 1558
rect 3570 1578 3630 1638
rect 3476 1538 3486 1552
rect 3426 1478 3486 1538
rect 3426 1438 3436 1478
rect 3476 1438 3486 1478
rect 3426 1422 3486 1438
rect 3570 1538 3580 1578
rect 3620 1538 3630 1578
rect 3570 1478 3630 1538
rect 3570 1438 3580 1478
rect 3620 1438 3630 1478
rect 3570 1422 3630 1438
rect 3858 1778 3918 1984
rect 3858 1738 3868 1778
rect 3908 1738 3918 1778
rect 3858 1678 3918 1738
rect 3858 1638 3868 1678
rect 3908 1638 3918 1678
rect 3858 1578 3918 1638
rect 4002 1778 4062 1828
rect 4002 1738 4012 1778
rect 4052 1738 4062 1778
rect 4002 1678 4062 1738
rect 4002 1638 4012 1678
rect 4052 1638 4062 1678
rect 4002 1616 4062 1638
rect 4146 1778 4206 1984
rect 4146 1738 4156 1778
rect 4196 1738 4206 1778
rect 4146 1678 4206 1738
rect 4146 1638 4156 1678
rect 4196 1638 4206 1678
rect 3858 1538 3868 1578
rect 3908 1538 3918 1578
rect 4000 1610 4064 1616
rect 4000 1558 4006 1610
rect 4058 1558 4064 1610
rect 4000 1552 4012 1558
rect 3858 1478 3918 1538
rect 3858 1438 3868 1478
rect 3908 1438 3918 1478
rect 3858 1422 3918 1438
rect 4002 1538 4012 1552
rect 4052 1552 4064 1558
rect 4146 1578 4206 1638
rect 4434 1778 4494 1828
rect 4434 1738 4444 1778
rect 4484 1738 4494 1778
rect 4578 1778 4638 1828
rect 4578 1760 4588 1778
rect 4434 1678 4494 1738
rect 4576 1754 4588 1760
rect 4628 1760 4638 1778
rect 4722 1778 4782 1828
rect 4628 1754 4640 1760
rect 4576 1702 4582 1754
rect 4634 1702 4640 1754
rect 4576 1696 4640 1702
rect 4722 1738 4732 1778
rect 4772 1738 4782 1778
rect 4434 1638 4444 1678
rect 4484 1638 4494 1678
rect 4434 1616 4494 1638
rect 4578 1678 4638 1696
rect 4578 1638 4588 1678
rect 4628 1638 4638 1678
rect 4052 1538 4062 1552
rect 4002 1478 4062 1538
rect 4002 1438 4012 1478
rect 4052 1438 4062 1478
rect 4002 1422 4062 1438
rect 4146 1538 4156 1578
rect 4196 1538 4206 1578
rect 4432 1610 4496 1616
rect 4432 1558 4438 1610
rect 4490 1558 4496 1610
rect 4432 1552 4444 1558
rect 4146 1478 4206 1538
rect 4146 1438 4156 1478
rect 4196 1438 4206 1478
rect 4146 1422 4206 1438
rect 4434 1538 4444 1552
rect 4484 1552 4496 1558
rect 4578 1578 4638 1638
rect 4722 1678 4782 1738
rect 4722 1638 4732 1678
rect 4772 1638 4782 1678
rect 4722 1616 4782 1638
rect 5010 1778 5070 1984
rect 5538 1982 5570 2044
rect 5664 1982 5708 2044
rect 5872 2042 5936 2048
rect 5872 1990 5878 2042
rect 5930 1990 5936 2042
rect 5872 1984 5936 1990
rect 6160 2042 6224 2048
rect 6160 1990 6166 2042
rect 6218 1990 6224 2042
rect 6160 1984 6224 1990
rect 5010 1738 5020 1778
rect 5060 1738 5070 1778
rect 5010 1678 5070 1738
rect 5010 1638 5020 1678
rect 5060 1638 5070 1678
rect 4484 1538 4494 1552
rect 4434 1478 4494 1538
rect 4434 1438 4444 1478
rect 4484 1438 4494 1478
rect 4434 1422 4494 1438
rect 4578 1538 4588 1578
rect 4628 1538 4638 1578
rect 4720 1610 4784 1616
rect 4720 1558 4726 1610
rect 4778 1558 4784 1610
rect 4720 1552 4732 1558
rect 4578 1478 4638 1538
rect 4578 1438 4588 1478
rect 4628 1438 4638 1478
rect 4578 1422 4638 1438
rect 4722 1538 4732 1552
rect 4772 1552 4784 1558
rect 5010 1578 5070 1638
rect 4772 1538 4782 1552
rect 4722 1478 4782 1538
rect 4722 1438 4732 1478
rect 4772 1438 4782 1478
rect 4722 1422 4782 1438
rect 5010 1538 5020 1578
rect 5060 1538 5070 1578
rect 5010 1478 5070 1538
rect 5010 1438 5020 1478
rect 5060 1438 5070 1478
rect 5010 1422 5070 1438
rect 5154 1778 5214 1828
rect 5154 1738 5164 1778
rect 5204 1738 5214 1778
rect 5298 1778 5358 1828
rect 5298 1760 5308 1778
rect 5154 1678 5214 1738
rect 5296 1754 5308 1760
rect 5348 1760 5358 1778
rect 5348 1754 5360 1760
rect 5296 1702 5302 1754
rect 5354 1702 5360 1754
rect 5296 1696 5360 1702
rect 5154 1638 5164 1678
rect 5204 1638 5214 1678
rect 5154 1578 5214 1638
rect 5154 1538 5164 1578
rect 5204 1538 5214 1578
rect 5154 1478 5214 1538
rect 5154 1438 5164 1478
rect 5204 1438 5214 1478
rect 5154 1422 5214 1438
rect 5298 1678 5358 1696
rect 5298 1638 5308 1678
rect 5348 1638 5358 1678
rect 5298 1578 5358 1638
rect 5298 1538 5308 1578
rect 5348 1538 5358 1578
rect 5298 1478 5358 1538
rect 5298 1438 5308 1478
rect 5348 1438 5358 1478
rect 5298 1422 5358 1438
rect 5538 1666 5708 1982
rect 5538 1476 5572 1666
rect 5652 1476 5708 1666
rect 5538 1424 5708 1476
rect 5874 1778 5934 1984
rect 5874 1738 5884 1778
rect 5924 1738 5934 1778
rect 5874 1678 5934 1738
rect 5874 1638 5884 1678
rect 5924 1638 5934 1678
rect 5874 1578 5934 1638
rect 6018 1778 6078 1828
rect 6018 1738 6028 1778
rect 6068 1738 6078 1778
rect 6018 1678 6078 1738
rect 6018 1638 6028 1678
rect 6068 1638 6078 1678
rect 6018 1616 6078 1638
rect 6162 1778 6222 1984
rect 6162 1738 6172 1778
rect 6212 1738 6222 1778
rect 6162 1678 6222 1738
rect 6162 1638 6172 1678
rect 6212 1638 6222 1678
rect 5874 1538 5884 1578
rect 5924 1538 5934 1578
rect 6016 1610 6080 1616
rect 6016 1558 6022 1610
rect 6074 1558 6080 1610
rect 6016 1552 6028 1558
rect 5874 1478 5934 1538
rect 5874 1438 5884 1478
rect 5924 1438 5934 1478
rect 5874 1422 5934 1438
rect 6018 1538 6028 1552
rect 6068 1552 6080 1558
rect 6162 1578 6222 1638
rect 6068 1538 6078 1552
rect 6018 1478 6078 1538
rect 6018 1438 6028 1478
rect 6068 1438 6078 1478
rect 6018 1422 6078 1438
rect 6162 1538 6172 1578
rect 6212 1538 6222 1578
rect 6162 1478 6222 1538
rect 6162 1438 6172 1478
rect 6212 1438 6222 1478
rect 6162 1422 6222 1438
rect 200 1322 374 1332
rect 200 1313 262 1322
rect 200 1279 220 1313
rect 254 1279 262 1313
rect 200 1270 262 1279
rect 314 1313 374 1322
rect 314 1279 328 1313
rect 362 1279 374 1313
rect 314 1270 374 1279
rect 200 1260 374 1270
rect 776 1322 950 1332
rect 776 1313 838 1322
rect 776 1279 796 1313
rect 830 1279 838 1313
rect 776 1270 838 1279
rect 890 1313 950 1322
rect 890 1279 904 1313
rect 938 1279 950 1313
rect 890 1270 950 1279
rect 776 1260 950 1270
rect 1352 1322 1526 1332
rect 1352 1313 1414 1322
rect 1352 1279 1372 1313
rect 1406 1279 1414 1313
rect 1352 1270 1414 1279
rect 1466 1313 1526 1322
rect 1466 1279 1480 1313
rect 1514 1279 1526 1313
rect 1466 1270 1526 1279
rect 1352 1260 1526 1270
rect 1928 1322 2102 1332
rect 1928 1313 1990 1322
rect 1928 1279 1948 1313
rect 1982 1279 1990 1313
rect 1928 1270 1990 1279
rect 2042 1313 2102 1322
rect 2042 1279 2056 1313
rect 2090 1279 2102 1313
rect 2042 1270 2102 1279
rect 1928 1260 2102 1270
rect 2414 1314 2504 1332
rect 2414 1278 2436 1314
rect 2472 1278 2504 1314
rect 2414 1260 2504 1278
rect 2678 1322 2768 1332
rect 2678 1270 2710 1322
rect 2762 1270 2768 1322
rect 2678 1260 2768 1270
rect 3368 1322 3542 1332
rect 3368 1313 3430 1322
rect 3368 1279 3388 1313
rect 3422 1279 3430 1313
rect 3368 1270 3430 1279
rect 3482 1313 3542 1322
rect 3482 1279 3496 1313
rect 3530 1279 3542 1313
rect 3482 1270 3542 1279
rect 3368 1260 3542 1270
rect 3944 1322 4118 1332
rect 3944 1313 4006 1322
rect 3944 1279 3964 1313
rect 3998 1279 4006 1313
rect 3944 1270 4006 1279
rect 4058 1313 4118 1322
rect 4058 1279 4072 1313
rect 4106 1279 4118 1313
rect 4058 1270 4118 1279
rect 3944 1260 4118 1270
rect 4520 1322 4694 1332
rect 4520 1313 4582 1322
rect 4520 1279 4540 1313
rect 4574 1279 4582 1313
rect 4520 1270 4582 1279
rect 4634 1313 4694 1322
rect 4634 1279 4648 1313
rect 4682 1279 4694 1313
rect 4634 1270 4694 1279
rect 4520 1260 4694 1270
rect 5006 1314 5096 1332
rect 5006 1278 5028 1314
rect 5064 1278 5096 1314
rect 5006 1260 5096 1278
rect 5270 1322 5360 1332
rect 5270 1270 5302 1322
rect 5354 1270 5360 1322
rect 5270 1260 5360 1270
rect 5960 1322 6134 1332
rect 5960 1313 6022 1322
rect 5960 1279 5980 1313
rect 6014 1279 6022 1313
rect 5960 1270 6022 1279
rect 6074 1313 6134 1322
rect 6074 1279 6088 1313
rect 6122 1279 6134 1313
rect 6074 1270 6134 1279
rect 5960 1260 6134 1270
rect 2418 1040 2478 1260
rect 5010 1040 5070 1260
rect 2416 1034 2480 1040
rect 2416 982 2422 1034
rect 2474 982 2480 1034
rect 2416 976 2480 982
rect 5008 1034 5072 1040
rect 5008 982 5014 1034
rect 5066 982 5072 1034
rect 5008 976 5072 982
rect 2418 756 2478 976
rect 5010 756 5070 976
rect 200 746 374 756
rect 200 737 262 746
rect 200 703 220 737
rect 254 703 262 737
rect 200 694 262 703
rect 314 737 374 746
rect 314 703 328 737
rect 362 703 374 737
rect 314 694 374 703
rect 200 684 374 694
rect 776 746 950 756
rect 776 737 838 746
rect 776 703 796 737
rect 830 703 838 737
rect 776 694 838 703
rect 890 737 950 746
rect 890 703 904 737
rect 938 703 950 737
rect 890 694 950 703
rect 776 684 950 694
rect 1352 746 1526 756
rect 1352 737 1414 746
rect 1352 703 1372 737
rect 1406 703 1414 737
rect 1352 694 1414 703
rect 1466 737 1526 746
rect 1466 703 1480 737
rect 1514 703 1526 737
rect 1466 694 1526 703
rect 1352 684 1526 694
rect 1928 746 2102 756
rect 1928 737 1990 746
rect 1928 703 1948 737
rect 1982 703 1990 737
rect 1928 694 1990 703
rect 2042 737 2102 746
rect 2042 703 2056 737
rect 2090 703 2102 737
rect 2042 694 2102 703
rect 1928 684 2102 694
rect 2414 738 2504 756
rect 2414 702 2436 738
rect 2472 702 2504 738
rect 2414 684 2504 702
rect 2678 746 2768 756
rect 2678 694 2710 746
rect 2762 694 2768 746
rect 2678 684 2768 694
rect 3368 746 3542 756
rect 3368 737 3430 746
rect 3368 703 3388 737
rect 3422 703 3430 737
rect 3368 694 3430 703
rect 3482 737 3542 746
rect 3482 703 3496 737
rect 3530 703 3542 737
rect 3482 694 3542 703
rect 3368 684 3542 694
rect 3944 746 4118 756
rect 3944 737 4006 746
rect 3944 703 3964 737
rect 3998 703 4006 737
rect 3944 694 4006 703
rect 4058 737 4118 746
rect 4058 703 4072 737
rect 4106 703 4118 737
rect 4058 694 4118 703
rect 3944 684 4118 694
rect 4520 746 4694 756
rect 4520 737 4582 746
rect 4520 703 4540 737
rect 4574 703 4582 737
rect 4520 694 4582 703
rect 4634 737 4694 746
rect 4634 703 4648 737
rect 4682 703 4694 737
rect 4634 694 4694 703
rect 4520 684 4694 694
rect 5006 738 5096 756
rect 5006 702 5028 738
rect 5064 702 5096 738
rect 5006 684 5096 702
rect 5270 746 5360 756
rect 5270 694 5302 746
rect 5354 694 5360 746
rect 5270 684 5360 694
rect 5960 746 6134 756
rect 5960 737 6022 746
rect 5960 703 5980 737
rect 6014 703 6022 737
rect 5960 694 6022 703
rect 6074 737 6134 746
rect 6074 703 6088 737
rect 6122 703 6134 737
rect 6074 694 6134 703
rect 5960 684 6134 694
rect 114 598 174 614
rect 114 558 124 598
rect 164 558 174 598
rect 114 498 174 558
rect 114 458 124 498
rect 164 458 174 498
rect 258 598 318 614
rect 258 558 268 598
rect 308 558 318 598
rect 258 498 318 558
rect 258 464 268 498
rect 114 32 174 458
rect 256 458 268 464
rect 308 464 318 498
rect 402 598 462 614
rect 402 558 412 598
rect 452 558 462 598
rect 402 498 462 558
rect 308 458 320 464
rect 256 406 262 458
rect 314 406 320 458
rect 256 400 320 406
rect 402 458 412 498
rect 452 458 462 498
rect 258 286 318 400
rect 402 32 462 458
rect 690 598 750 614
rect 690 558 700 598
rect 740 558 750 598
rect 690 498 750 558
rect 690 458 700 498
rect 740 458 750 498
rect 834 598 894 614
rect 834 558 844 598
rect 884 558 894 598
rect 834 498 894 558
rect 834 464 844 498
rect 690 32 750 458
rect 832 458 844 464
rect 884 464 894 498
rect 978 598 1038 614
rect 978 558 988 598
rect 1028 558 1038 598
rect 978 498 1038 558
rect 884 458 896 464
rect 832 406 838 458
rect 890 406 896 458
rect 832 400 896 406
rect 978 458 988 498
rect 1028 458 1038 498
rect 834 286 894 400
rect 978 32 1038 458
rect 1266 598 1326 614
rect 1266 558 1276 598
rect 1316 558 1326 598
rect 1266 498 1326 558
rect 1266 458 1276 498
rect 1316 458 1326 498
rect 1410 598 1470 614
rect 1410 558 1420 598
rect 1460 558 1470 598
rect 1410 498 1470 558
rect 1410 464 1420 498
rect 1266 32 1326 458
rect 1408 458 1420 464
rect 1460 464 1470 498
rect 1554 598 1614 614
rect 1554 558 1564 598
rect 1604 558 1614 598
rect 1554 498 1614 558
rect 1460 458 1472 464
rect 1408 406 1414 458
rect 1466 406 1472 458
rect 1408 400 1472 406
rect 1554 458 1564 498
rect 1604 458 1614 498
rect 1842 598 1902 614
rect 1842 558 1852 598
rect 1892 558 1902 598
rect 1842 498 1902 558
rect 1842 464 1852 498
rect 1410 286 1470 400
rect 1554 32 1614 458
rect 1840 458 1852 464
rect 1892 464 1902 498
rect 1986 598 2046 614
rect 1986 558 1996 598
rect 2036 558 2046 598
rect 1986 498 2046 558
rect 1892 458 1904 464
rect 1840 406 1846 458
rect 1898 406 1904 458
rect 1840 400 1904 406
rect 1986 458 1996 498
rect 2036 458 2046 498
rect 2130 598 2190 614
rect 2130 558 2140 598
rect 2180 558 2190 598
rect 2130 498 2190 558
rect 2130 464 2140 498
rect 1842 286 1902 400
rect 1986 320 2046 458
rect 2128 458 2140 464
rect 2180 464 2190 498
rect 2418 598 2478 614
rect 2418 558 2428 598
rect 2468 558 2478 598
rect 2418 498 2478 558
rect 2180 458 2192 464
rect 2128 406 2134 458
rect 2186 406 2192 458
rect 2128 400 2192 406
rect 2418 458 2428 498
rect 2468 458 2478 498
rect 1984 314 2048 320
rect 1984 262 1990 314
rect 2042 262 2048 314
rect 2130 286 2190 400
rect 1984 256 2048 262
rect 2418 32 2478 458
rect 2562 598 2622 614
rect 2562 558 2572 598
rect 2612 558 2622 598
rect 2562 498 2622 558
rect 2562 458 2572 498
rect 2612 458 2622 498
rect 2562 442 2622 458
rect 2706 598 2766 614
rect 2706 558 2716 598
rect 2756 558 2766 598
rect 2706 498 2766 558
rect 2706 458 2716 498
rect 2756 458 2766 498
rect 2706 320 2766 458
rect 3282 598 3342 614
rect 3282 558 3292 598
rect 3332 558 3342 598
rect 3282 498 3342 558
rect 3282 458 3292 498
rect 3332 458 3342 498
rect 3426 598 3486 614
rect 3426 558 3436 598
rect 3476 558 3486 598
rect 3426 498 3486 558
rect 3426 464 3436 498
rect 2704 314 2768 320
rect 2704 262 2710 314
rect 2762 262 2768 314
rect 2704 256 2768 262
rect 3282 32 3342 458
rect 3424 458 3436 464
rect 3476 464 3486 498
rect 3570 598 3630 614
rect 3570 558 3580 598
rect 3620 558 3630 598
rect 3570 498 3630 558
rect 3476 458 3488 464
rect 3424 406 3430 458
rect 3482 406 3488 458
rect 3424 400 3488 406
rect 3570 458 3580 498
rect 3620 458 3630 498
rect 3426 286 3486 400
rect 3570 32 3630 458
rect 3858 598 3918 614
rect 3858 558 3868 598
rect 3908 558 3918 598
rect 3858 498 3918 558
rect 3858 458 3868 498
rect 3908 458 3918 498
rect 4002 598 4062 614
rect 4002 558 4012 598
rect 4052 558 4062 598
rect 4002 498 4062 558
rect 4002 464 4012 498
rect 3858 32 3918 458
rect 4000 458 4012 464
rect 4052 464 4062 498
rect 4146 598 4206 614
rect 4146 558 4156 598
rect 4196 558 4206 598
rect 4146 498 4206 558
rect 4052 458 4064 464
rect 4000 406 4006 458
rect 4058 406 4064 458
rect 4000 400 4064 406
rect 4146 458 4156 498
rect 4196 458 4206 498
rect 4434 598 4494 614
rect 4434 558 4444 598
rect 4484 558 4494 598
rect 4434 498 4494 558
rect 4434 464 4444 498
rect 4002 286 4062 400
rect 4146 32 4206 458
rect 4432 458 4444 464
rect 4484 464 4494 498
rect 4578 598 4638 614
rect 4578 558 4588 598
rect 4628 558 4638 598
rect 4578 498 4638 558
rect 4484 458 4496 464
rect 4432 406 4438 458
rect 4490 406 4496 458
rect 4432 400 4496 406
rect 4578 458 4588 498
rect 4628 458 4638 498
rect 4722 598 4782 614
rect 4722 558 4732 598
rect 4772 558 4782 598
rect 4722 498 4782 558
rect 4722 464 4732 498
rect 4434 286 4494 400
rect 4578 320 4638 458
rect 4720 458 4732 464
rect 4772 464 4782 498
rect 5010 598 5070 614
rect 5010 558 5020 598
rect 5060 558 5070 598
rect 5010 498 5070 558
rect 4772 458 4784 464
rect 4720 406 4726 458
rect 4778 406 4784 458
rect 4720 400 4784 406
rect 5010 458 5020 498
rect 5060 458 5070 498
rect 4576 314 4640 320
rect 4576 262 4582 314
rect 4634 262 4640 314
rect 4722 286 4782 400
rect 4576 256 4640 262
rect 5010 32 5070 458
rect 5154 598 5214 614
rect 5154 558 5164 598
rect 5204 558 5214 598
rect 5154 498 5214 558
rect 5154 458 5164 498
rect 5204 458 5214 498
rect 5154 442 5214 458
rect 5298 598 5358 614
rect 5298 558 5308 598
rect 5348 558 5358 598
rect 5298 498 5358 558
rect 5298 458 5308 498
rect 5348 458 5358 498
rect 5298 320 5358 458
rect 5542 592 5756 642
rect 5542 450 5600 592
rect 5710 450 5756 592
rect 5296 314 5360 320
rect 5296 262 5302 314
rect 5354 262 5360 314
rect 5296 256 5360 262
rect 5542 40 5756 450
rect 112 26 176 32
rect 112 -26 118 26
rect 170 -26 176 26
rect 112 -32 176 -26
rect 400 26 464 32
rect 400 -26 406 26
rect 458 -26 464 26
rect 400 -32 464 -26
rect 688 26 752 32
rect 688 -26 694 26
rect 746 -26 752 26
rect 688 -32 752 -26
rect 976 26 1040 32
rect 976 -26 982 26
rect 1034 -26 1040 26
rect 976 -32 1040 -26
rect 1264 26 1328 32
rect 1264 -26 1270 26
rect 1322 -26 1328 26
rect 1264 -32 1328 -26
rect 1552 26 1616 32
rect 1552 -26 1558 26
rect 1610 -26 1616 26
rect 1552 -32 1616 -26
rect 2416 26 2480 32
rect 2416 -26 2422 26
rect 2474 -26 2480 26
rect 2416 -32 2480 -26
rect 3280 26 3344 32
rect 3280 -26 3286 26
rect 3338 -26 3344 26
rect 3280 -32 3344 -26
rect 3568 26 3632 32
rect 3568 -26 3574 26
rect 3626 -26 3632 26
rect 3568 -32 3632 -26
rect 3856 26 3920 32
rect 3856 -26 3862 26
rect 3914 -26 3920 26
rect 3856 -32 3920 -26
rect 4144 26 4208 32
rect 4144 -26 4150 26
rect 4202 -26 4208 26
rect 4144 -32 4208 -26
rect 5008 26 5072 32
rect 5008 -26 5014 26
rect 5066 -26 5072 26
rect 5008 -32 5072 -26
rect 114 -40 174 -32
rect 402 -40 462 -32
rect 690 -40 750 -32
rect 978 -40 1038 -32
rect 1266 -40 1326 -32
rect 1554 -40 1614 -32
rect 3282 -40 3342 -32
rect 3570 -40 3630 -32
rect 3858 -40 3918 -32
rect 4146 -40 4206 -32
rect 5542 -38 5604 40
rect 5702 -38 5756 40
rect 5874 598 5934 614
rect 5874 558 5884 598
rect 5924 558 5934 598
rect 5874 498 5934 558
rect 5874 458 5884 498
rect 5924 458 5934 498
rect 6018 598 6078 614
rect 6018 558 6028 598
rect 6068 558 6078 598
rect 6018 498 6078 558
rect 6018 464 6028 498
rect 5874 32 5934 458
rect 6016 458 6028 464
rect 6068 464 6078 498
rect 6162 598 6222 614
rect 6162 558 6172 598
rect 6212 558 6222 598
rect 6162 498 6222 558
rect 6068 458 6080 464
rect 6016 406 6022 458
rect 6074 406 6080 458
rect 6016 400 6080 406
rect 6162 458 6172 498
rect 6212 458 6222 498
rect 6018 286 6078 400
rect 6162 32 6222 458
rect 5872 26 5936 32
rect 5872 -26 5878 26
rect 5930 -26 5936 26
rect 5872 -32 5936 -26
rect 6160 26 6224 32
rect 6160 -26 6166 26
rect 6218 -26 6224 26
rect 6160 -32 6224 -26
rect 5874 -40 5934 -32
rect 6162 -40 6222 -32
<< via1 >>
rect 118 1990 170 2042
rect 406 1990 458 2042
rect 694 1990 746 2042
rect 982 1990 1034 2042
rect 1270 1990 1322 2042
rect 1558 1990 1610 2042
rect 2422 1990 2474 2042
rect 3286 1990 3338 2042
rect 3574 1990 3626 2042
rect 3862 1990 3914 2042
rect 4150 1990 4202 2042
rect 5014 1990 5066 2042
rect 262 1578 314 1610
rect 262 1558 268 1578
rect 268 1558 308 1578
rect 308 1558 314 1578
rect 838 1578 890 1610
rect 838 1558 844 1578
rect 844 1558 884 1578
rect 884 1558 890 1578
rect 1414 1578 1466 1610
rect 1414 1558 1420 1578
rect 1420 1558 1460 1578
rect 1460 1558 1466 1578
rect 1990 1738 1996 1754
rect 1996 1738 2036 1754
rect 2036 1738 2042 1754
rect 1990 1702 2042 1738
rect 1846 1578 1898 1610
rect 1846 1558 1852 1578
rect 1852 1558 1892 1578
rect 1892 1558 1898 1578
rect 2134 1578 2186 1610
rect 2134 1558 2140 1578
rect 2140 1558 2180 1578
rect 2180 1558 2186 1578
rect 2710 1738 2716 1754
rect 2716 1738 2756 1754
rect 2756 1738 2762 1754
rect 2710 1702 2762 1738
rect 3430 1578 3482 1610
rect 3430 1558 3436 1578
rect 3436 1558 3476 1578
rect 3476 1558 3482 1578
rect 4006 1578 4058 1610
rect 4006 1558 4012 1578
rect 4012 1558 4052 1578
rect 4052 1558 4058 1578
rect 4582 1738 4588 1754
rect 4588 1738 4628 1754
rect 4628 1738 4634 1754
rect 4582 1702 4634 1738
rect 4438 1578 4490 1610
rect 4438 1558 4444 1578
rect 4444 1558 4484 1578
rect 4484 1558 4490 1578
rect 5570 1982 5664 2044
rect 5878 1990 5930 2042
rect 6166 1990 6218 2042
rect 4726 1578 4778 1610
rect 4726 1558 4732 1578
rect 4732 1558 4772 1578
rect 4772 1558 4778 1578
rect 5302 1738 5308 1754
rect 5308 1738 5348 1754
rect 5348 1738 5354 1754
rect 5302 1702 5354 1738
rect 6022 1578 6074 1610
rect 6022 1558 6028 1578
rect 6028 1558 6068 1578
rect 6068 1558 6074 1578
rect 262 1270 314 1322
rect 838 1270 890 1322
rect 1414 1270 1466 1322
rect 1990 1270 2042 1322
rect 2710 1314 2762 1322
rect 2710 1278 2720 1314
rect 2720 1278 2756 1314
rect 2756 1278 2762 1314
rect 2710 1270 2762 1278
rect 3430 1270 3482 1322
rect 4006 1270 4058 1322
rect 4582 1270 4634 1322
rect 5302 1314 5354 1322
rect 5302 1278 5312 1314
rect 5312 1278 5348 1314
rect 5348 1278 5354 1314
rect 5302 1270 5354 1278
rect 6022 1270 6074 1322
rect 2422 982 2474 1034
rect 5014 982 5066 1034
rect 262 694 314 746
rect 838 694 890 746
rect 1414 694 1466 746
rect 1990 694 2042 746
rect 2710 738 2762 746
rect 2710 702 2714 738
rect 2714 702 2750 738
rect 2750 702 2762 738
rect 2710 694 2762 702
rect 3430 694 3482 746
rect 4006 694 4058 746
rect 4582 694 4634 746
rect 5302 738 5354 746
rect 5302 702 5306 738
rect 5306 702 5342 738
rect 5342 702 5354 738
rect 5302 694 5354 702
rect 6022 694 6074 746
rect 262 406 314 458
rect 838 406 890 458
rect 1414 406 1466 458
rect 1846 406 1898 458
rect 2134 406 2186 458
rect 1990 262 2042 314
rect 2710 262 2762 314
rect 3430 406 3482 458
rect 4006 406 4058 458
rect 4438 406 4490 458
rect 4726 406 4778 458
rect 4582 262 4634 314
rect 5302 262 5354 314
rect 118 -26 170 26
rect 406 -26 458 26
rect 694 -26 746 26
rect 982 -26 1034 26
rect 1270 -26 1322 26
rect 1558 -26 1610 26
rect 2422 -26 2474 26
rect 3286 -26 3338 26
rect 3574 -26 3626 26
rect 3862 -26 3914 26
rect 4150 -26 4202 26
rect 5014 -26 5066 26
rect 5604 -38 5702 40
rect 6022 406 6074 458
rect 5878 -26 5930 26
rect 6166 -26 6218 26
<< metal2 >>
rect -40 2044 6376 2076
rect -40 2042 5570 2044
rect -40 1990 118 2042
rect 170 1990 406 2042
rect 458 1990 694 2042
rect 746 1990 982 2042
rect 1034 1990 1270 2042
rect 1322 1990 1558 2042
rect 1610 1990 2422 2042
rect 2474 1990 3286 2042
rect 3338 1990 3574 2042
rect 3626 1990 3862 2042
rect 3914 1990 4150 2042
rect 4202 1990 5014 2042
rect 5066 1990 5570 2042
rect -40 1982 5570 1990
rect 5664 2042 6376 2044
rect 5664 1990 5878 2042
rect 5930 1990 6166 2042
rect 6218 1990 6376 2042
rect 5664 1982 6376 1990
rect -40 1956 6376 1982
rect 1978 1758 2054 1766
rect 1836 1756 2196 1758
rect 1836 1700 1988 1756
rect 2044 1700 2196 1756
rect 1836 1698 2196 1700
rect 2698 1756 2774 1766
rect 4570 1758 4646 1766
rect 2698 1700 2708 1756
rect 2764 1700 2774 1756
rect 1978 1690 2054 1698
rect 2698 1690 2774 1700
rect 4428 1756 4788 1758
rect 4428 1700 4580 1756
rect 4636 1700 4788 1756
rect 4428 1698 4788 1700
rect 5290 1756 5366 1766
rect 5290 1700 5300 1756
rect 5356 1700 5366 1756
rect 4570 1690 4646 1698
rect 5290 1690 5366 1700
rect 250 1614 326 1622
rect 826 1614 902 1622
rect 1408 1614 1472 1616
rect 1840 1614 1904 1616
rect 2128 1614 2192 1616
rect 3418 1614 3494 1622
rect 4000 1614 4064 1616
rect 4432 1614 4496 1616
rect 4720 1614 4784 1616
rect 6010 1614 6086 1622
rect 108 1612 468 1614
rect 108 1556 260 1612
rect 316 1556 468 1612
rect 108 1554 468 1556
rect 684 1612 1044 1614
rect 684 1556 836 1612
rect 892 1556 1044 1612
rect 684 1554 1044 1556
rect 1260 1610 2236 1614
rect 1260 1558 1414 1610
rect 1466 1558 1846 1610
rect 1898 1558 2134 1610
rect 2186 1558 2236 1610
rect 1260 1554 2236 1558
rect 3276 1612 3636 1614
rect 3276 1556 3428 1612
rect 3484 1556 3636 1612
rect 3276 1554 3636 1556
rect 3852 1610 4828 1614
rect 3852 1558 4006 1610
rect 4058 1558 4438 1610
rect 4490 1558 4726 1610
rect 4778 1558 4828 1610
rect 3852 1554 4828 1558
rect 5868 1612 6228 1614
rect 5868 1556 6020 1612
rect 6076 1556 6228 1612
rect 5868 1554 6228 1556
rect 250 1546 326 1554
rect 826 1546 902 1554
rect 1408 1552 1472 1554
rect 1840 1552 1904 1554
rect 2128 1552 2192 1554
rect 3418 1546 3494 1554
rect 4000 1552 4064 1554
rect 4432 1552 4496 1554
rect 4720 1552 4784 1554
rect 6010 1546 6086 1554
rect 106 1326 182 1334
rect 256 1326 320 1328
rect 682 1326 758 1334
rect 832 1326 896 1328
rect 1402 1326 1478 1334
rect 1834 1326 1910 1334
rect 1984 1326 2048 1328
rect 2554 1326 2630 1334
rect 2704 1326 2768 1328
rect 106 1324 468 1326
rect 106 1268 116 1324
rect 172 1322 468 1324
rect 172 1270 262 1322
rect 314 1270 468 1322
rect 172 1268 468 1270
rect 106 1266 468 1268
rect 682 1324 1044 1326
rect 682 1268 692 1324
rect 748 1322 1044 1324
rect 748 1270 838 1322
rect 890 1270 1044 1322
rect 748 1268 1044 1270
rect 682 1266 1044 1268
rect 1260 1324 1620 1326
rect 1260 1268 1412 1324
rect 1468 1268 1620 1324
rect 1260 1266 1620 1268
rect 1834 1324 2196 1326
rect 1834 1268 1844 1324
rect 1900 1322 2196 1324
rect 1900 1270 1990 1322
rect 2042 1270 2196 1322
rect 1900 1268 2196 1270
rect 1834 1266 2196 1268
rect 2554 1324 2768 1326
rect 2554 1268 2564 1324
rect 2620 1322 2768 1324
rect 2620 1270 2710 1322
rect 2762 1270 2768 1322
rect 2620 1268 2768 1270
rect 2554 1266 2768 1268
rect 106 1258 182 1266
rect 256 1264 320 1266
rect 682 1258 758 1266
rect 832 1264 896 1266
rect 1402 1258 1478 1266
rect 1834 1258 1910 1266
rect 1984 1264 2048 1266
rect 2554 1258 2630 1266
rect 2704 1264 2768 1266
rect 3274 1326 3350 1334
rect 3424 1326 3488 1328
rect 3994 1326 4070 1334
rect 4426 1326 4502 1334
rect 4576 1326 4640 1328
rect 5146 1326 5222 1334
rect 5296 1326 5360 1328
rect 3274 1324 3636 1326
rect 3274 1268 3284 1324
rect 3340 1322 3636 1324
rect 3340 1270 3430 1322
rect 3482 1270 3636 1322
rect 3340 1268 3636 1270
rect 3274 1266 3636 1268
rect 3852 1324 4212 1326
rect 3852 1268 4004 1324
rect 4060 1268 4212 1324
rect 3852 1266 4212 1268
rect 4426 1324 4788 1326
rect 4426 1268 4436 1324
rect 4492 1322 4788 1324
rect 4492 1270 4582 1322
rect 4634 1270 4788 1322
rect 4492 1268 4788 1270
rect 4426 1266 4788 1268
rect 5146 1324 5360 1326
rect 5146 1268 5156 1324
rect 5212 1322 5360 1324
rect 5212 1270 5302 1322
rect 5354 1270 5360 1322
rect 5212 1268 5360 1270
rect 5146 1266 5360 1268
rect 3274 1258 3350 1266
rect 3424 1264 3488 1266
rect 3994 1258 4070 1266
rect 4426 1258 4502 1266
rect 4576 1264 4640 1266
rect 5146 1258 5222 1266
rect 5296 1264 5360 1266
rect 5866 1326 5942 1334
rect 6016 1326 6080 1328
rect 5866 1324 6228 1326
rect 5866 1268 5876 1324
rect 5932 1322 6228 1324
rect 5932 1270 6022 1322
rect 6074 1270 6228 1322
rect 5932 1268 6228 1270
rect 5866 1266 6228 1268
rect 5866 1258 5942 1266
rect 6016 1264 6080 1266
rect 2410 1038 2486 1046
rect 5002 1038 5078 1046
rect 2410 1036 2756 1038
rect 2410 980 2420 1036
rect 2476 980 2756 1036
rect 2410 978 2756 980
rect 5002 1036 5348 1038
rect 5002 980 5012 1036
rect 5068 980 5348 1036
rect 5002 978 5348 980
rect 2410 970 2486 978
rect 5002 970 5078 978
rect 106 750 182 758
rect 256 750 320 752
rect 682 750 758 758
rect 832 750 896 752
rect 1402 750 1478 758
rect 1984 750 2048 752
rect 2122 750 2198 758
rect 106 748 468 750
rect 106 692 116 748
rect 172 746 468 748
rect 172 694 262 746
rect 314 694 468 746
rect 172 692 468 694
rect 106 690 468 692
rect 682 748 1044 750
rect 682 692 692 748
rect 748 746 1044 748
rect 748 694 838 746
rect 890 694 1044 746
rect 748 692 1044 694
rect 682 690 1044 692
rect 1260 748 1620 750
rect 1260 692 1412 748
rect 1468 692 1620 748
rect 1260 690 1620 692
rect 1836 748 2198 750
rect 1836 746 2132 748
rect 1836 694 1990 746
rect 2042 694 2132 746
rect 1836 692 2132 694
rect 2188 692 2198 748
rect 1836 690 2198 692
rect 106 682 182 690
rect 256 688 320 690
rect 682 682 758 690
rect 832 688 896 690
rect 1402 682 1478 690
rect 1984 688 2048 690
rect 2122 682 2198 690
rect 2704 750 2768 752
rect 2842 750 2918 758
rect 2704 748 2918 750
rect 2704 746 2852 748
rect 2704 694 2710 746
rect 2762 694 2852 746
rect 2704 692 2852 694
rect 2908 692 2918 748
rect 2704 690 2918 692
rect 2704 688 2768 690
rect 2842 682 2918 690
rect 3274 750 3350 758
rect 3424 750 3488 752
rect 3994 750 4070 758
rect 4576 750 4640 752
rect 4714 750 4790 758
rect 3274 748 3636 750
rect 3274 692 3284 748
rect 3340 746 3636 748
rect 3340 694 3430 746
rect 3482 694 3636 746
rect 3340 692 3636 694
rect 3274 690 3636 692
rect 3852 748 4212 750
rect 3852 692 4004 748
rect 4060 692 4212 748
rect 3852 690 4212 692
rect 4428 748 4790 750
rect 4428 746 4724 748
rect 4428 694 4582 746
rect 4634 694 4724 746
rect 4428 692 4724 694
rect 4780 692 4790 748
rect 4428 690 4790 692
rect 3274 682 3350 690
rect 3424 688 3488 690
rect 3994 682 4070 690
rect 4576 688 4640 690
rect 4714 682 4790 690
rect 5296 750 5360 752
rect 5434 750 5510 758
rect 5296 748 5510 750
rect 5296 746 5444 748
rect 5296 694 5302 746
rect 5354 694 5444 746
rect 5296 692 5444 694
rect 5500 692 5510 748
rect 5296 690 5510 692
rect 5296 688 5360 690
rect 5434 682 5510 690
rect 5866 750 5942 758
rect 6016 750 6080 752
rect 5866 748 6228 750
rect 5866 692 5876 748
rect 5932 746 6228 748
rect 5932 694 6022 746
rect 6074 694 6228 746
rect 5932 692 6228 694
rect 5866 690 6228 692
rect 5866 682 5942 690
rect 6016 688 6080 690
rect 250 462 326 470
rect 826 462 902 470
rect 1408 462 1472 464
rect 1840 462 1904 464
rect 2128 462 2192 464
rect 3418 462 3494 470
rect 4000 462 4064 464
rect 4432 462 4496 464
rect 4720 462 4784 464
rect 6010 462 6086 470
rect 108 460 468 462
rect 108 404 260 460
rect 316 404 468 460
rect 108 402 468 404
rect 684 460 1044 462
rect 684 404 836 460
rect 892 404 1044 460
rect 684 402 1044 404
rect 1260 458 2236 462
rect 1260 406 1414 458
rect 1466 406 1846 458
rect 1898 406 2134 458
rect 2186 406 2236 458
rect 1260 402 2236 406
rect 3276 460 3636 462
rect 3276 404 3428 460
rect 3484 404 3636 460
rect 3276 402 3636 404
rect 3852 458 4828 462
rect 3852 406 4006 458
rect 4058 406 4438 458
rect 4490 406 4726 458
rect 4778 406 4828 458
rect 3852 402 4828 406
rect 5868 460 6228 462
rect 5868 404 6020 460
rect 6076 404 6228 460
rect 5868 402 6228 404
rect 250 394 326 402
rect 826 394 902 402
rect 1408 400 1472 402
rect 1840 400 1904 402
rect 2128 400 2192 402
rect 3418 394 3494 402
rect 4000 400 4064 402
rect 4432 400 4496 402
rect 4720 400 4784 402
rect 6010 394 6086 402
rect 1978 318 2054 326
rect 1836 316 2196 318
rect 1836 260 1988 316
rect 2044 260 2196 316
rect 1836 258 2196 260
rect 2698 316 2774 326
rect 4570 318 4646 326
rect 2698 260 2708 316
rect 2764 260 2774 316
rect 1978 250 2054 258
rect 2698 250 2774 260
rect 4428 316 4788 318
rect 4428 260 4580 316
rect 4636 260 4788 316
rect 4428 258 4788 260
rect 5290 316 5366 326
rect 5290 260 5300 316
rect 5356 260 5366 316
rect 4570 250 4646 258
rect 5290 250 5366 260
rect -40 40 6376 60
rect -40 26 5604 40
rect -40 -26 118 26
rect 170 -26 406 26
rect 458 -26 694 26
rect 746 -26 982 26
rect 1034 -26 1270 26
rect 1322 -26 1558 26
rect 1610 -26 2422 26
rect 2474 -26 3286 26
rect 3338 -26 3574 26
rect 3626 -26 3862 26
rect 3914 -26 4150 26
rect 4202 -26 5014 26
rect 5066 -26 5604 26
rect -40 -38 5604 -26
rect 5702 26 6376 40
rect 5702 -26 5878 26
rect 5930 -26 6166 26
rect 6218 -26 6376 26
rect 5702 -38 6376 -26
rect -40 -60 6376 -38
<< via2 >>
rect 1988 1754 2044 1756
rect 1988 1702 1990 1754
rect 1990 1702 2042 1754
rect 2042 1702 2044 1754
rect 1988 1700 2044 1702
rect 2708 1754 2764 1756
rect 2708 1702 2710 1754
rect 2710 1702 2762 1754
rect 2762 1702 2764 1754
rect 2708 1700 2764 1702
rect 4580 1754 4636 1756
rect 4580 1702 4582 1754
rect 4582 1702 4634 1754
rect 4634 1702 4636 1754
rect 4580 1700 4636 1702
rect 5300 1754 5356 1756
rect 5300 1702 5302 1754
rect 5302 1702 5354 1754
rect 5354 1702 5356 1754
rect 5300 1700 5356 1702
rect 260 1610 316 1612
rect 260 1558 262 1610
rect 262 1558 314 1610
rect 314 1558 316 1610
rect 260 1556 316 1558
rect 836 1610 892 1612
rect 836 1558 838 1610
rect 838 1558 890 1610
rect 890 1558 892 1610
rect 836 1556 892 1558
rect 3428 1610 3484 1612
rect 3428 1558 3430 1610
rect 3430 1558 3482 1610
rect 3482 1558 3484 1610
rect 3428 1556 3484 1558
rect 6020 1610 6076 1612
rect 6020 1558 6022 1610
rect 6022 1558 6074 1610
rect 6074 1558 6076 1610
rect 6020 1556 6076 1558
rect 116 1268 172 1324
rect 692 1268 748 1324
rect 1412 1322 1468 1324
rect 1412 1270 1414 1322
rect 1414 1270 1466 1322
rect 1466 1270 1468 1322
rect 1412 1268 1468 1270
rect 1844 1268 1900 1324
rect 2564 1268 2620 1324
rect 3284 1268 3340 1324
rect 4004 1322 4060 1324
rect 4004 1270 4006 1322
rect 4006 1270 4058 1322
rect 4058 1270 4060 1322
rect 4004 1268 4060 1270
rect 4436 1268 4492 1324
rect 5156 1268 5212 1324
rect 5876 1268 5932 1324
rect 2420 1034 2476 1036
rect 2420 982 2422 1034
rect 2422 982 2474 1034
rect 2474 982 2476 1034
rect 2420 980 2476 982
rect 5012 1034 5068 1036
rect 5012 982 5014 1034
rect 5014 982 5066 1034
rect 5066 982 5068 1034
rect 5012 980 5068 982
rect 116 692 172 748
rect 692 692 748 748
rect 1412 746 1468 748
rect 1412 694 1414 746
rect 1414 694 1466 746
rect 1466 694 1468 746
rect 1412 692 1468 694
rect 2132 692 2188 748
rect 2852 692 2908 748
rect 3284 692 3340 748
rect 4004 746 4060 748
rect 4004 694 4006 746
rect 4006 694 4058 746
rect 4058 694 4060 746
rect 4004 692 4060 694
rect 4724 692 4780 748
rect 5444 692 5500 748
rect 5876 692 5932 748
rect 260 458 316 460
rect 260 406 262 458
rect 262 406 314 458
rect 314 406 316 458
rect 260 404 316 406
rect 836 458 892 460
rect 836 406 838 458
rect 838 406 890 458
rect 890 406 892 458
rect 836 404 892 406
rect 3428 458 3484 460
rect 3428 406 3430 458
rect 3430 406 3482 458
rect 3482 406 3484 458
rect 3428 404 3484 406
rect 6020 458 6076 460
rect 6020 406 6022 458
rect 6022 406 6074 458
rect 6074 406 6076 458
rect 6020 404 6076 406
rect 1988 314 2044 316
rect 1988 262 1990 314
rect 1990 262 2042 314
rect 2042 262 2044 314
rect 1988 260 2044 262
rect 2708 314 2764 316
rect 2708 262 2710 314
rect 2710 262 2762 314
rect 2762 262 2764 314
rect 2708 260 2764 262
rect 4580 314 4636 316
rect 4580 262 4582 314
rect 4582 262 4634 314
rect 4634 262 4636 314
rect 4580 260 4636 262
rect 5300 314 5356 316
rect 5300 262 5302 314
rect 5302 262 5354 314
rect 5354 262 5356 314
rect 5300 260 5356 262
<< metal3 >>
rect 1978 1756 2054 1766
rect 1978 1700 1988 1756
rect 2044 1700 2054 1756
rect 1978 1690 2054 1700
rect 2698 1756 2774 1766
rect 2698 1700 2708 1756
rect 2764 1700 2774 1756
rect 2698 1690 2774 1700
rect 4570 1756 4646 1766
rect 4570 1700 4580 1756
rect 4636 1700 4646 1756
rect 4570 1690 4646 1700
rect 5290 1756 5366 1766
rect 5290 1700 5300 1756
rect 5356 1700 5366 1756
rect 5290 1690 5366 1700
rect 250 1612 326 1622
rect 250 1556 260 1612
rect 316 1556 326 1612
rect 250 1546 326 1556
rect 826 1612 902 1622
rect 826 1556 836 1612
rect 892 1556 902 1612
rect 826 1546 902 1556
rect 106 1324 182 1334
rect 106 1268 116 1324
rect 172 1268 182 1324
rect 106 1258 182 1268
rect 114 758 174 1258
rect 106 748 182 758
rect 106 692 116 748
rect 172 692 182 748
rect 106 682 182 692
rect 258 470 318 1546
rect 682 1324 758 1334
rect 682 1268 692 1324
rect 748 1268 758 1324
rect 682 1258 758 1268
rect 690 758 750 1258
rect 682 748 758 758
rect 682 692 692 748
rect 748 692 758 748
rect 682 682 758 692
rect 250 460 326 470
rect 250 404 260 460
rect 316 404 326 460
rect 250 394 326 404
rect 258 326 318 394
rect 690 326 750 682
rect 834 470 894 1546
rect 1402 1324 1478 1334
rect 1402 1268 1412 1324
rect 1468 1268 1478 1324
rect 1402 1258 1478 1268
rect 1834 1324 1910 1334
rect 1834 1268 1844 1324
rect 1900 1268 1910 1324
rect 1834 1258 1910 1268
rect 1410 758 1470 1258
rect 1402 748 1478 758
rect 1402 692 1412 748
rect 1468 692 1478 748
rect 1402 682 1478 692
rect 826 460 902 470
rect 826 404 836 460
rect 892 404 902 460
rect 826 394 902 404
rect 250 320 326 326
rect 250 256 256 320
rect 320 256 326 320
rect 250 250 326 256
rect 682 320 758 326
rect 682 256 688 320
rect 752 256 758 320
rect 682 250 758 256
rect 834 182 894 394
rect 1842 182 1902 1258
rect 1986 470 2046 1690
rect 2130 758 2190 1326
rect 2418 1046 2478 1326
rect 2554 1324 2630 1334
rect 2554 1268 2564 1324
rect 2620 1268 2630 1324
rect 2554 1258 2630 1268
rect 2410 1036 2486 1046
rect 2410 980 2420 1036
rect 2476 980 2486 1036
rect 2410 970 2486 980
rect 2122 748 2198 758
rect 2122 692 2132 748
rect 2188 692 2198 748
rect 2122 682 2198 692
rect 1978 464 2054 470
rect 1978 400 1984 464
rect 2048 400 2054 464
rect 1978 394 2054 400
rect 1986 326 2046 394
rect 2130 326 2190 682
rect 2418 614 2478 970
rect 2410 608 2486 614
rect 2410 544 2416 608
rect 2480 544 2486 608
rect 2410 538 2486 544
rect 2562 326 2622 1258
rect 2706 470 2766 1690
rect 3418 1612 3494 1622
rect 3418 1556 3428 1612
rect 3484 1556 3494 1612
rect 3418 1546 3494 1556
rect 2850 758 2910 1326
rect 3274 1324 3350 1334
rect 3274 1268 3284 1324
rect 3340 1268 3350 1324
rect 3274 1258 3350 1268
rect 3282 758 3342 1258
rect 2842 748 2918 758
rect 2842 692 2852 748
rect 2908 692 2918 748
rect 2842 682 2918 692
rect 3274 748 3350 758
rect 3274 692 3284 748
rect 3340 692 3350 748
rect 3274 682 3350 692
rect 2698 464 2774 470
rect 2698 400 2704 464
rect 2768 400 2774 464
rect 2698 394 2774 400
rect 2706 326 2766 394
rect 1978 316 2054 326
rect 1978 260 1988 316
rect 2044 260 2054 316
rect 1978 250 2054 260
rect 2122 320 2198 326
rect 2122 256 2128 320
rect 2192 256 2198 320
rect 2122 250 2198 256
rect 2554 320 2630 326
rect 2554 256 2560 320
rect 2624 256 2630 320
rect 2554 250 2630 256
rect 2698 316 2774 326
rect 2698 260 2708 316
rect 2764 260 2774 316
rect 2698 250 2774 260
rect 2850 182 2910 682
rect 3282 470 3342 682
rect 3426 614 3486 1546
rect 3994 1324 4070 1334
rect 3994 1268 4004 1324
rect 4060 1268 4070 1324
rect 3994 1258 4070 1268
rect 4426 1324 4502 1334
rect 4426 1268 4436 1324
rect 4492 1268 4502 1324
rect 4426 1258 4502 1268
rect 4002 758 4062 1258
rect 3994 748 4070 758
rect 3994 692 4004 748
rect 4060 692 4070 748
rect 3994 682 4070 692
rect 4002 614 4062 682
rect 3418 608 3494 614
rect 3418 544 3424 608
rect 3488 544 3494 608
rect 3418 538 3494 544
rect 3994 608 4070 614
rect 3994 544 4000 608
rect 4064 544 4070 608
rect 3994 538 4070 544
rect 3426 470 3486 538
rect 3274 464 3350 470
rect 3274 400 3280 464
rect 3344 400 3350 464
rect 3274 394 3350 400
rect 3418 460 3494 470
rect 3418 404 3428 460
rect 3484 404 3494 460
rect 3418 394 3494 404
rect 4434 326 4494 1258
rect 4578 470 4638 1690
rect 4722 758 4782 1326
rect 5010 1046 5070 1326
rect 5146 1324 5222 1334
rect 5146 1268 5156 1324
rect 5212 1268 5222 1324
rect 5146 1258 5222 1268
rect 5002 1036 5078 1046
rect 5002 980 5012 1036
rect 5068 980 5078 1036
rect 5002 970 5078 980
rect 4714 748 4790 758
rect 4714 692 4724 748
rect 4780 692 4790 748
rect 4714 682 4790 692
rect 4570 464 4646 470
rect 4570 400 4576 464
rect 4640 400 4646 464
rect 4570 394 4646 400
rect 4578 326 4638 394
rect 4426 320 4502 326
rect 4426 256 4432 320
rect 4496 256 4502 320
rect 4426 250 4502 256
rect 4570 316 4646 326
rect 4570 260 4580 316
rect 4636 260 4646 316
rect 4570 250 4646 260
rect 4722 182 4782 682
rect 5010 614 5070 970
rect 5002 608 5078 614
rect 5002 544 5008 608
rect 5072 544 5078 608
rect 5002 538 5078 544
rect 5154 182 5214 1258
rect 5298 470 5358 1690
rect 6010 1612 6086 1622
rect 6010 1556 6020 1612
rect 6076 1556 6086 1612
rect 6010 1546 6086 1556
rect 5442 758 5502 1326
rect 5866 1324 5942 1334
rect 5866 1268 5876 1324
rect 5932 1268 5942 1324
rect 5866 1258 5942 1268
rect 5874 758 5934 1258
rect 5434 748 5510 758
rect 5434 692 5444 748
rect 5500 692 5510 748
rect 5434 682 5510 692
rect 5866 748 5942 758
rect 5866 692 5876 748
rect 5932 692 5942 748
rect 5866 682 5942 692
rect 5290 464 5366 470
rect 5290 400 5296 464
rect 5360 400 5366 464
rect 5290 394 5366 400
rect 5298 326 5358 394
rect 5442 326 5502 682
rect 5874 470 5934 682
rect 6018 614 6078 1546
rect 6010 608 6086 614
rect 6010 544 6016 608
rect 6080 544 6086 608
rect 6010 538 6086 544
rect 6018 470 6078 538
rect 5866 464 5942 470
rect 5866 400 5872 464
rect 5936 400 5942 464
rect 5866 394 5942 400
rect 6010 460 6086 470
rect 6010 404 6020 460
rect 6076 404 6086 460
rect 6010 394 6086 404
rect 5290 316 5366 326
rect 5290 260 5300 316
rect 5356 260 5366 316
rect 5290 250 5366 260
rect 5434 320 5510 326
rect 5434 256 5440 320
rect 5504 256 5510 320
rect 5434 250 5510 256
rect 826 176 902 182
rect 826 112 832 176
rect 896 112 902 176
rect 826 106 902 112
rect 1834 176 1910 182
rect 1834 112 1840 176
rect 1904 112 1910 176
rect 1834 106 1910 112
rect 2842 176 2918 182
rect 2842 112 2848 176
rect 2912 112 2918 176
rect 2842 106 2918 112
rect 4714 176 4790 182
rect 4714 112 4720 176
rect 4784 112 4790 176
rect 4714 106 4790 112
rect 5146 176 5222 182
rect 5146 112 5152 176
rect 5216 112 5222 176
rect 5146 106 5222 112
<< via3 >>
rect 256 256 320 320
rect 688 256 752 320
rect 1984 400 2048 464
rect 2416 544 2480 608
rect 2704 400 2768 464
rect 2128 256 2192 320
rect 2560 256 2624 320
rect 3424 544 3488 608
rect 4000 544 4064 608
rect 3280 400 3344 464
rect 4576 400 4640 464
rect 4432 256 4496 320
rect 5008 544 5072 608
rect 5296 400 5360 464
rect 6016 544 6080 608
rect 5872 400 5936 464
rect 5440 256 5504 320
rect 832 112 896 176
rect 1840 112 1904 176
rect 2848 112 2912 176
rect 4720 112 4784 176
rect 5152 112 5216 176
<< metal4 >>
rect 2414 608 2482 610
rect 2414 544 2416 608
rect 2480 606 2482 608
rect 3422 608 3490 610
rect 3422 606 3424 608
rect 2480 546 3424 606
rect 2480 544 2482 546
rect 2414 542 2482 544
rect 3422 544 3424 546
rect 3488 606 3490 608
rect 3998 608 4066 610
rect 3998 606 4000 608
rect 3488 546 4000 606
rect 3488 544 3490 546
rect 3422 542 3490 544
rect 3998 544 4000 546
rect 4064 544 4066 608
rect 3998 542 4066 544
rect 5006 608 5074 610
rect 5006 544 5008 608
rect 5072 606 5074 608
rect 6014 608 6082 610
rect 6014 606 6016 608
rect 5072 546 6016 606
rect 5072 544 5074 546
rect 5006 542 5074 544
rect 6014 544 6016 546
rect 6080 544 6082 608
rect 6014 542 6082 544
rect 1982 464 2050 466
rect 1982 400 1984 464
rect 2048 462 2050 464
rect 2702 464 2770 466
rect 2702 462 2704 464
rect 2048 402 2704 462
rect 2048 400 2050 402
rect 1982 398 2050 400
rect 2702 400 2704 402
rect 2768 462 2770 464
rect 3278 464 3346 466
rect 3278 462 3280 464
rect 2768 402 3280 462
rect 2768 400 2770 402
rect 2702 398 2770 400
rect 3278 400 3280 402
rect 3344 400 3346 464
rect 3278 398 3346 400
rect 4574 464 4642 466
rect 4574 400 4576 464
rect 4640 462 4642 464
rect 5294 464 5362 466
rect 5294 462 5296 464
rect 4640 402 5296 462
rect 4640 400 4642 402
rect 4574 398 4642 400
rect 5294 400 5296 402
rect 5360 462 5362 464
rect 5870 464 5938 466
rect 5870 462 5872 464
rect 5360 402 5872 462
rect 5360 400 5362 402
rect 5294 398 5362 400
rect 5870 400 5872 402
rect 5936 400 5938 464
rect 5870 398 5938 400
rect 254 320 322 322
rect 254 256 256 320
rect 320 318 322 320
rect 686 320 754 322
rect 686 318 688 320
rect 320 258 688 318
rect 320 256 322 258
rect 254 254 322 256
rect 686 256 688 258
rect 752 318 754 320
rect 2126 320 2194 322
rect 2126 318 2128 320
rect 752 258 2128 318
rect 752 256 754 258
rect 686 254 754 256
rect 2126 256 2128 258
rect 2192 318 2194 320
rect 2558 320 2626 322
rect 2558 318 2560 320
rect 2192 258 2560 318
rect 2192 256 2194 258
rect 2126 254 2194 256
rect 2558 256 2560 258
rect 2624 318 2626 320
rect 4430 320 4498 322
rect 4430 318 4432 320
rect 2624 258 4432 318
rect 2624 256 2626 258
rect 2558 254 2626 256
rect 4430 256 4432 258
rect 4496 318 4498 320
rect 5438 320 5506 322
rect 5438 318 5440 320
rect 4496 258 5440 318
rect 4496 256 4498 258
rect 4430 254 4498 256
rect 5438 256 5440 258
rect 5504 256 5506 320
rect 5438 254 5506 256
rect 830 176 898 178
rect 830 112 832 176
rect 896 174 898 176
rect 1838 176 1906 178
rect 1838 174 1840 176
rect 896 114 1840 174
rect 896 112 898 114
rect 830 110 898 112
rect 1838 112 1840 114
rect 1904 174 1906 176
rect 2846 176 2914 178
rect 2846 174 2848 176
rect 1904 114 2848 174
rect 1904 112 1906 114
rect 1838 110 1906 112
rect 2846 112 2848 114
rect 2912 174 2914 176
rect 4718 176 4786 178
rect 4718 174 4720 176
rect 2912 114 4720 174
rect 2912 112 2914 114
rect 2846 110 2914 112
rect 4718 112 4720 114
rect 4784 174 4786 176
rect 5150 176 5218 178
rect 5150 174 5152 176
rect 4784 114 5152 174
rect 4784 112 4786 114
rect 4718 110 4786 112
rect 5150 112 5152 114
rect 5216 112 5218 176
rect 5150 110 5218 112
<< labels >>
flabel metal3 1440 1008 1440 1008 0 FreeSans 480 90 0 0 I
flabel metal3 144 1008 144 1008 0 FreeSans 480 90 0 0 CLK
flabel metal3 6048 1008 6048 1008 0 FreeSans 480 90 0 0 O
flabel metal2 3168 0 3168 0 0 FreeSans 960 0 0 0 VSS
flabel metal2 3168 2016 3168 2016 0 FreeSans 960 0 0 0 VDD
flabel metal3 144 1008 144 1008 0 FreeSans 480 90 0 0 inv0/I
flabel metal3 288 1008 288 1008 0 FreeSans 480 90 0 0 inv0/O
flabel metal2 288 0 288 0 0 FreeSans 960 0 0 0 inv0/VSS
flabel metal2 288 2016 288 2016 0 FreeSans 960 0 0 0 inv0/VDD
flabel space 0 0 144 1008 0 FreeSans 320 90 0 0 inv0/MN0_IBNDL0/nmos_boundary
flabel space 432 0 576 1008 0 FreeSans 320 90 0 0 inv0/MN0_IBNDR0/nmos_boundary
flabel metal1 114 288 174 614 0 FreeSans 240 0 0 0 inv0/MN0_IM0/S0
flabel metal1 258 288 318 614 0 FreeSans 240 0 0 0 inv0/MN0_IM0/D0
flabel metal1 402 288 462 614 0 FreeSans 240 0 0 0 inv0/MN0_IM0/S1
flabel metal1 200 684 374 756 0 FreeSans 240 0 0 0 inv0/MN0_IM0/G0
rlabel pwell 104 654 134 676 1 inv0/MN0_IM0/BODY
flabel space 0 1008 144 2016 0 FreeSans 320 90 0 0 inv0/MP0_IBNDL0/pmos_boundary
flabel space 432 1008 576 2016 0 FreeSans 320 90 0 0 inv0/MP0_IBNDR0/pmos_boundary
flabel metal1 258 1422 318 1828 0 FreeSans 160 0 0 0 inv0/MP0_IM0/D0
flabel metal1 200 1260 374 1332 0 FreeSans 160 0 0 0 inv0/MP0_IM0/G0
flabel metal1 114 1422 174 1828 0 FreeSans 160 0 0 0 inv0/MP0_IM0/S0
flabel metal1 402 1422 462 1828 0 FreeSans 160 0 0 0 inv0/MP0_IM0/S1
flabel nwell 124 1346 148 1362 0 FreeSans 80 0 0 0 inv0/MP0_IM0/BODY
flabel metal3 720 1008 720 1008 0 FreeSans 480 90 0 0 inv1/I
flabel metal3 864 1008 864 1008 0 FreeSans 480 90 0 0 inv1/O
flabel metal2 864 0 864 0 0 FreeSans 960 0 0 0 inv1/VSS
flabel metal2 864 2016 864 2016 0 FreeSans 960 0 0 0 inv1/VDD
flabel space 576 0 720 1008 0 FreeSans 320 90 0 0 inv1/MN0_IBNDL0/nmos_boundary
flabel space 1008 0 1152 1008 0 FreeSans 320 90 0 0 inv1/MN0_IBNDR0/nmos_boundary
flabel metal1 690 288 750 614 0 FreeSans 240 0 0 0 inv1/MN0_IM0/S0
flabel metal1 834 288 894 614 0 FreeSans 240 0 0 0 inv1/MN0_IM0/D0
flabel metal1 978 288 1038 614 0 FreeSans 240 0 0 0 inv1/MN0_IM0/S1
flabel metal1 776 684 950 756 0 FreeSans 240 0 0 0 inv1/MN0_IM0/G0
rlabel pwell 680 654 710 676 1 inv1/MN0_IM0/BODY
flabel space 576 1008 720 2016 0 FreeSans 320 90 0 0 inv1/MP0_IBNDL0/pmos_boundary
flabel space 1008 1008 1152 2016 0 FreeSans 320 90 0 0 inv1/MP0_IBNDR0/pmos_boundary
flabel metal1 834 1422 894 1828 0 FreeSans 160 0 0 0 inv1/MP0_IM0/D0
flabel metal1 776 1260 950 1332 0 FreeSans 160 0 0 0 inv1/MP0_IM0/G0
flabel metal1 690 1422 750 1828 0 FreeSans 160 0 0 0 inv1/MP0_IM0/S0
flabel metal1 978 1422 1038 1828 0 FreeSans 160 0 0 0 inv1/MP0_IM0/S1
flabel nwell 700 1346 724 1362 0 FreeSans 80 0 0 0 inv1/MP0_IM0/BODY
flabel metal3 1440 1008 1440 1008 0 FreeSans 480 90 0 0 tinv0/I
flabel metal3 2160 1008 2160 1008 0 FreeSans 480 90 0 0 tinv0/EN
flabel metal3 1872 1008 1872 1008 0 FreeSans 480 90 0 0 tinv0/ENB
flabel metal3 2016 1008 2016 1008 0 FreeSans 480 90 0 0 tinv0/O
flabel metal2 1728 0 1728 0 0 FreeSans 960 0 0 0 tinv0/VSS
flabel metal2 1728 2016 1728 2016 0 FreeSans 960 0 0 0 tinv0/VDD
flabel space 1152 0 1296 1008 0 FreeSans 320 90 0 0 tinv0/MN0_IBNDL0/nmos_boundary
flabel space 1584 0 1728 1008 0 FreeSans 320 90 0 0 tinv0/MN0_IBNDR0/nmos_boundary
flabel metal1 1266 288 1326 614 0 FreeSans 240 0 0 0 tinv0/MN0_IM0/S0
flabel metal1 1410 288 1470 614 0 FreeSans 240 0 0 0 tinv0/MN0_IM0/D0
flabel metal1 1554 288 1614 614 0 FreeSans 240 0 0 0 tinv0/MN0_IM0/S1
flabel metal1 1352 684 1526 756 0 FreeSans 240 0 0 0 tinv0/MN0_IM0/G0
rlabel pwell 1256 654 1286 676 1 tinv0/MN0_IM0/BODY
flabel space 1728 0 1872 1008 0 FreeSans 320 90 0 0 tinv0/MN1_IBNDL0/nmos_boundary
flabel metal1 1842 288 1902 614 0 FreeSans 240 0 0 0 tinv0/MN1_IM0/S0
flabel metal1 1986 288 2046 614 0 FreeSans 240 0 0 0 tinv0/MN1_IM0/D0
flabel metal1 2130 288 2190 614 0 FreeSans 240 0 0 0 tinv0/MN1_IM0/S1
flabel metal1 1928 684 2102 756 0 FreeSans 240 0 0 0 tinv0/MN1_IM0/G0
rlabel pwell 1832 654 1862 676 1 tinv0/MN1_IM0/BODY
flabel space 2160 0 2304 1008 0 FreeSans 320 90 0 0 tinv0/MN1_IBNDR0/nmos_boundary
flabel space 1152 1008 1296 2016 0 FreeSans 320 90 0 0 tinv0/MP0_IBNDL0/pmos_boundary
flabel space 1584 1008 1728 2016 0 FreeSans 320 90 0 0 tinv0/MP0_IBNDR0/pmos_boundary
flabel metal1 1410 1422 1470 1828 0 FreeSans 160 0 0 0 tinv0/MP0_IM0/D0
flabel metal1 1352 1260 1526 1332 0 FreeSans 160 0 0 0 tinv0/MP0_IM0/G0
flabel metal1 1266 1422 1326 1828 0 FreeSans 160 0 0 0 tinv0/MP0_IM0/S0
flabel metal1 1554 1422 1614 1828 0 FreeSans 160 0 0 0 tinv0/MP0_IM0/S1
flabel nwell 1276 1346 1300 1362 0 FreeSans 80 0 0 0 tinv0/MP0_IM0/BODY
flabel space 1728 1008 1872 2016 0 FreeSans 320 90 0 0 tinv0/MP1_IBNDL0/pmos_boundary
flabel metal1 1986 1422 2046 1828 0 FreeSans 160 0 0 0 tinv0/MP1_IM0/D0
flabel metal1 1928 1260 2102 1332 0 FreeSans 160 0 0 0 tinv0/MP1_IM0/G0
flabel metal1 1842 1422 1902 1828 0 FreeSans 160 0 0 0 tinv0/MP1_IM0/S0
flabel metal1 2130 1422 2190 1828 0 FreeSans 160 0 0 0 tinv0/MP1_IM0/S1
flabel nwell 1852 1346 1876 1362 0 FreeSans 80 0 0 0 tinv0/MP1_IM0/BODY
flabel space 2160 1008 2304 2016 0 FreeSans 320 90 0 0 tinv0/MP1_IBNDR0/pmos_boundary
flabel metal3 2448 1008 2448 1008 0 FreeSans 480 90 0 0 tinv_small0/I
flabel metal3 2736 1008 2736 1008 0 FreeSans 480 90 0 0 tinv_small0/O
flabel metal3 2880 1008 2880 1008 0 FreeSans 480 90 0 0 tinv_small0/EN
flabel metal3 2592 1008 2592 1008 0 FreeSans 480 90 0 0 tinv_small0/ENB
flabel metal2 2736 0 2736 0 0 FreeSans 960 0 0 0 tinv_small0/VSS
flabel metal2 2736 2016 2736 2016 0 FreeSans 960 0 0 0 tinv_small0/VDD
flabel space 2736 0 2880 1008 0 FreeSans 320 90 0 0 tinv_small0/nbndr/nmos_boundary
flabel space 2304 0 2448 1008 0 FreeSans 320 90 0 0 tinv_small0/nbndl/nmos_boundary
flabel space 3024 0 3168 1008 0 FreeSans 320 90 0 0 tinv_small0/nspace1/NMOS_SPACE
flabel space 2880 0 3024 1008 0 FreeSans 320 90 0 0 tinv_small0/nspace0/NMOS_SPACE
flabel metal1 2414 684 2504 756 0 FreeSans 160 0 0 0 tinv_small0/nstack/G0
flabel metal1 2678 684 2768 756 0 FreeSans 160 0 0 0 tinv_small0/nstack/G1
flabel metal1 2418 288 2478 614 0 FreeSans 160 0 0 0 tinv_small0/nstack/S0
rlabel pwell 2408 654 2438 676 1 tinv_small0/nstack/BODY
flabel metal1 2706 288 2766 614 0 FreeSans 160 0 0 0 tinv_small0/nstack/D0
flabel space 2736 1008 2880 2016 0 FreeSans 320 90 0 0 tinv_small0/pbndr/pmos_boundary
flabel space 2304 1008 2448 2016 0 FreeSans 320 90 0 0 tinv_small0/pbndl/pmos_boundary
flabel space 3024 1008 3168 2016 0 FreeSans 320 90 0 0 tinv_small0/pspace1/PMOS_SPACE
flabel space 2880 1008 3024 2016 0 FreeSans 320 90 0 0 tinv_small0/pspace0/PMOS_SPACE
flabel metal1 2414 1260 2504 1332 0 FreeSans 160 0 0 0 tinv_small0/pstack/G0
flabel metal1 2678 1260 2768 1332 0 FreeSans 160 0 0 0 tinv_small0/pstack/G1
flabel metal1 2418 1422 2478 1828 0 FreeSans 160 0 0 0 tinv_small0/pstack/S0
flabel nwell 2428 1346 2452 1362 0 FreeSans 80 0 0 0 tinv_small0/pstack/BODY
flabel metal1 2706 1422 2766 1828 0 FreeSans 160 0 0 0 tinv_small0/pstack/D0
flabel metal3 3312 1008 3312 1008 0 FreeSans 480 90 0 0 inv2/I
flabel metal3 3456 1008 3456 1008 0 FreeSans 480 90 0 0 inv2/O
flabel metal2 3456 0 3456 0 0 FreeSans 960 0 0 0 inv2/VSS
flabel metal2 3456 2016 3456 2016 0 FreeSans 960 0 0 0 inv2/VDD
flabel space 3168 0 3312 1008 0 FreeSans 320 90 0 0 inv2/MN0_IBNDL0/nmos_boundary
flabel space 3600 0 3744 1008 0 FreeSans 320 90 0 0 inv2/MN0_IBNDR0/nmos_boundary
flabel metal1 3282 288 3342 614 0 FreeSans 240 0 0 0 inv2/MN0_IM0/S0
flabel metal1 3426 288 3486 614 0 FreeSans 240 0 0 0 inv2/MN0_IM0/D0
flabel metal1 3570 288 3630 614 0 FreeSans 240 0 0 0 inv2/MN0_IM0/S1
flabel metal1 3368 684 3542 756 0 FreeSans 240 0 0 0 inv2/MN0_IM0/G0
rlabel pwell 3272 654 3302 676 1 inv2/MN0_IM0/BODY
flabel space 3168 1008 3312 2016 0 FreeSans 320 90 0 0 inv2/MP0_IBNDL0/pmos_boundary
flabel space 3600 1008 3744 2016 0 FreeSans 320 90 0 0 inv2/MP0_IBNDR0/pmos_boundary
flabel metal1 3426 1422 3486 1828 0 FreeSans 160 0 0 0 inv2/MP0_IM0/D0
flabel metal1 3368 1260 3542 1332 0 FreeSans 160 0 0 0 inv2/MP0_IM0/G0
flabel metal1 3282 1422 3342 1828 0 FreeSans 160 0 0 0 inv2/MP0_IM0/S0
flabel metal1 3570 1422 3630 1828 0 FreeSans 160 0 0 0 inv2/MP0_IM0/S1
flabel nwell 3292 1346 3316 1362 0 FreeSans 80 0 0 0 inv2/MP0_IM0/BODY
flabel metal3 4032 1008 4032 1008 0 FreeSans 480 90 0 0 tinv1/I
flabel metal3 4752 1008 4752 1008 0 FreeSans 480 90 0 0 tinv1/EN
flabel metal3 4464 1008 4464 1008 0 FreeSans 480 90 0 0 tinv1/ENB
flabel metal3 4608 1008 4608 1008 0 FreeSans 480 90 0 0 tinv1/O
flabel metal2 4320 0 4320 0 0 FreeSans 960 0 0 0 tinv1/VSS
flabel metal2 4320 2016 4320 2016 0 FreeSans 960 0 0 0 tinv1/VDD
flabel space 3744 0 3888 1008 0 FreeSans 320 90 0 0 tinv1/MN0_IBNDL0/nmos_boundary
flabel space 4176 0 4320 1008 0 FreeSans 320 90 0 0 tinv1/MN0_IBNDR0/nmos_boundary
flabel metal1 3858 288 3918 614 0 FreeSans 240 0 0 0 tinv1/MN0_IM0/S0
flabel metal1 4002 288 4062 614 0 FreeSans 240 0 0 0 tinv1/MN0_IM0/D0
flabel metal1 4146 288 4206 614 0 FreeSans 240 0 0 0 tinv1/MN0_IM0/S1
flabel metal1 3944 684 4118 756 0 FreeSans 240 0 0 0 tinv1/MN0_IM0/G0
rlabel pwell 3848 654 3878 676 1 tinv1/MN0_IM0/BODY
flabel space 4320 0 4464 1008 0 FreeSans 320 90 0 0 tinv1/MN1_IBNDL0/nmos_boundary
flabel metal1 4434 288 4494 614 0 FreeSans 240 0 0 0 tinv1/MN1_IM0/S0
flabel metal1 4578 288 4638 614 0 FreeSans 240 0 0 0 tinv1/MN1_IM0/D0
flabel metal1 4722 288 4782 614 0 FreeSans 240 0 0 0 tinv1/MN1_IM0/S1
flabel metal1 4520 684 4694 756 0 FreeSans 240 0 0 0 tinv1/MN1_IM0/G0
rlabel pwell 4424 654 4454 676 1 tinv1/MN1_IM0/BODY
flabel space 4752 0 4896 1008 0 FreeSans 320 90 0 0 tinv1/MN1_IBNDR0/nmos_boundary
flabel space 3744 1008 3888 2016 0 FreeSans 320 90 0 0 tinv1/MP0_IBNDL0/pmos_boundary
flabel space 4176 1008 4320 2016 0 FreeSans 320 90 0 0 tinv1/MP0_IBNDR0/pmos_boundary
flabel metal1 4002 1422 4062 1828 0 FreeSans 160 0 0 0 tinv1/MP0_IM0/D0
flabel metal1 3944 1260 4118 1332 0 FreeSans 160 0 0 0 tinv1/MP0_IM0/G0
flabel metal1 3858 1422 3918 1828 0 FreeSans 160 0 0 0 tinv1/MP0_IM0/S0
flabel metal1 4146 1422 4206 1828 0 FreeSans 160 0 0 0 tinv1/MP0_IM0/S1
flabel nwell 3868 1346 3892 1362 0 FreeSans 80 0 0 0 tinv1/MP0_IM0/BODY
flabel space 4320 1008 4464 2016 0 FreeSans 320 90 0 0 tinv1/MP1_IBNDL0/pmos_boundary
flabel metal1 4578 1422 4638 1828 0 FreeSans 160 0 0 0 tinv1/MP1_IM0/D0
flabel metal1 4520 1260 4694 1332 0 FreeSans 160 0 0 0 tinv1/MP1_IM0/G0
flabel metal1 4434 1422 4494 1828 0 FreeSans 160 0 0 0 tinv1/MP1_IM0/S0
flabel metal1 4722 1422 4782 1828 0 FreeSans 160 0 0 0 tinv1/MP1_IM0/S1
flabel nwell 4444 1346 4468 1362 0 FreeSans 80 0 0 0 tinv1/MP1_IM0/BODY
flabel space 4752 1008 4896 2016 0 FreeSans 320 90 0 0 tinv1/MP1_IBNDR0/pmos_boundary
flabel metal3 5040 1008 5040 1008 0 FreeSans 480 90 0 0 tinv_small1/I
flabel metal3 5328 1008 5328 1008 0 FreeSans 480 90 0 0 tinv_small1/O
flabel metal3 5472 1008 5472 1008 0 FreeSans 480 90 0 0 tinv_small1/EN
flabel metal3 5184 1008 5184 1008 0 FreeSans 480 90 0 0 tinv_small1/ENB
flabel metal2 5328 0 5328 0 0 FreeSans 960 0 0 0 tinv_small1/VSS
flabel metal2 5328 2016 5328 2016 0 FreeSans 960 0 0 0 tinv_small1/VDD
flabel space 5328 0 5472 1008 0 FreeSans 320 90 0 0 tinv_small1/nbndr/nmos_boundary
flabel space 4896 0 5040 1008 0 FreeSans 320 90 0 0 tinv_small1/nbndl/nmos_boundary
flabel space 5616 0 5760 1008 0 FreeSans 320 90 0 0 tinv_small1/nspace1/NMOS_SPACE
flabel space 5472 0 5616 1008 0 FreeSans 320 90 0 0 tinv_small1/nspace0/NMOS_SPACE
flabel metal1 5006 684 5096 756 0 FreeSans 160 0 0 0 tinv_small1/nstack/G0
flabel metal1 5270 684 5360 756 0 FreeSans 160 0 0 0 tinv_small1/nstack/G1
flabel metal1 5010 288 5070 614 0 FreeSans 160 0 0 0 tinv_small1/nstack/S0
rlabel pwell 5000 654 5030 676 1 tinv_small1/nstack/BODY
flabel metal1 5298 288 5358 614 0 FreeSans 160 0 0 0 tinv_small1/nstack/D0
flabel space 5328 1008 5472 2016 0 FreeSans 320 90 0 0 tinv_small1/pbndr/pmos_boundary
flabel space 4896 1008 5040 2016 0 FreeSans 320 90 0 0 tinv_small1/pbndl/pmos_boundary
flabel space 5616 1008 5760 2016 0 FreeSans 320 90 0 0 tinv_small1/pspace1/PMOS_SPACE
flabel space 5472 1008 5616 2016 0 FreeSans 320 90 0 0 tinv_small1/pspace0/PMOS_SPACE
flabel metal1 5006 1260 5096 1332 0 FreeSans 160 0 0 0 tinv_small1/pstack/G0
flabel metal1 5270 1260 5360 1332 0 FreeSans 160 0 0 0 tinv_small1/pstack/G1
flabel metal1 5010 1422 5070 1828 0 FreeSans 160 0 0 0 tinv_small1/pstack/S0
flabel nwell 5020 1346 5044 1362 0 FreeSans 80 0 0 0 tinv_small1/pstack/BODY
flabel metal1 5298 1422 5358 1828 0 FreeSans 160 0 0 0 tinv_small1/pstack/D0
flabel metal3 5904 1008 5904 1008 0 FreeSans 480 90 0 0 inv3/I
flabel metal3 6048 1008 6048 1008 0 FreeSans 480 90 0 0 inv3/O
flabel metal2 6048 0 6048 0 0 FreeSans 960 0 0 0 inv3/VSS
flabel metal2 6048 2016 6048 2016 0 FreeSans 960 0 0 0 inv3/VDD
flabel space 5760 0 5904 1008 0 FreeSans 320 90 0 0 inv3/MN0_IBNDL0/nmos_boundary
flabel space 6192 0 6336 1008 0 FreeSans 320 90 0 0 inv3/MN0_IBNDR0/nmos_boundary
flabel metal1 5874 288 5934 614 0 FreeSans 240 0 0 0 inv3/MN0_IM0/S0
flabel metal1 6018 288 6078 614 0 FreeSans 240 0 0 0 inv3/MN0_IM0/D0
flabel metal1 6162 288 6222 614 0 FreeSans 240 0 0 0 inv3/MN0_IM0/S1
flabel metal1 5960 684 6134 756 0 FreeSans 240 0 0 0 inv3/MN0_IM0/G0
rlabel pwell 5864 654 5894 676 1 inv3/MN0_IM0/BODY
flabel space 5760 1008 5904 2016 0 FreeSans 320 90 0 0 inv3/MP0_IBNDL0/pmos_boundary
flabel space 6192 1008 6336 2016 0 FreeSans 320 90 0 0 inv3/MP0_IBNDR0/pmos_boundary
flabel metal1 6018 1422 6078 1828 0 FreeSans 160 0 0 0 inv3/MP0_IM0/D0
flabel metal1 5960 1260 6134 1332 0 FreeSans 160 0 0 0 inv3/MP0_IM0/G0
flabel metal1 5874 1422 5934 1828 0 FreeSans 160 0 0 0 inv3/MP0_IM0/S0
flabel metal1 6162 1422 6222 1828 0 FreeSans 160 0 0 0 inv3/MP0_IM0/S1
flabel nwell 5884 1346 5908 1362 0 FreeSans 80 0 0 0 inv3/MP0_IM0/BODY
<< end >>
