magic
tech sky130A
magscale 1 2
timestamp 1706182685
<< error_p >>
rect -37 28 37 34
rect -37 -28 -28 28
rect -37 -34 37 -28
<< metal2 >>
rect -37 -28 -28 28
rect 28 -28 37 28
<< via2 >>
rect -28 -28 28 28
<< metal3 >>
rect -37 28 37 34
rect -37 -28 -28 28
rect 28 -28 37 28
rect -37 -34 37 -28
<< end >>
