magic
tech sky130A
timestamp 1655825056
<< pwell >>
rect 0 186 144 342
<< labels >>
flabel space 0 0 144 504 0 FreeSans 160 90 0 0 NMOS_SPACE_2X
<< end >>
