magic
tech sky130A
magscale 1 2
timestamp 1647160568
<< pwell >>
rect -56 304 224 440
<< nmoslvt >>
rect 26 330 56 414
rect 112 330 142 414
<< ndiff >>
rect -30 395 26 414
rect -30 361 -19 395
rect 15 361 26 395
rect -30 330 26 361
rect 56 395 112 414
rect 56 361 67 395
rect 101 361 112 395
rect 56 330 112 361
rect 142 395 198 414
rect 142 361 153 395
rect 187 361 198 395
rect 142 330 198 361
<< ndiffc >>
rect -19 361 15 395
rect 67 361 101 395
rect 153 361 187 395
<< poly >>
rect 17 495 151 511
rect 17 461 33 495
rect 67 461 101 495
rect 135 461 151 495
rect 17 445 151 461
rect 26 440 142 445
rect 26 414 56 440
rect 112 414 142 440
rect 26 304 56 330
rect 112 304 142 330
<< polycont >>
rect 33 461 67 495
rect 101 461 135 495
<< locali >>
rect 17 495 151 511
rect 17 461 31 495
rect 67 461 101 495
rect 137 461 151 495
rect 17 445 151 461
rect -19 395 15 411
rect -19 345 15 361
rect 67 395 101 411
rect 67 345 101 361
rect 153 395 187 411
rect 153 345 187 361
<< viali >>
rect 31 461 33 495
rect 33 461 65 495
rect 103 461 135 495
rect 135 461 137 495
rect -19 361 15 395
rect 67 361 101 395
rect 153 361 187 395
<< metal1 >>
rect 19 495 149 507
rect 19 461 31 495
rect 65 461 103 495
rect 137 461 149 495
rect 19 449 149 461
rect -25 395 21 414
rect -25 361 -19 395
rect 15 361 21 395
rect -25 265 21 361
rect 58 408 110 414
rect 58 345 110 356
rect 147 395 193 414
rect 147 361 153 395
rect 187 361 193 395
rect 147 265 193 361
rect -25 205 193 265
<< via1 >>
rect 58 395 110 408
rect 58 361 67 395
rect 67 361 101 395
rect 101 361 110 395
rect 58 356 110 361
<< metal2 >>
rect 58 408 110 414
rect 58 345 110 356
<< end >>
