magic
tech sky130A
magscale 1 2
timestamp 1708415439
<< checkpaint >>
rect -1260 2117 1704 2156
rect -1277 -799 1704 2117
rect -1277 -1289 1645 -799
rect -1260 -1344 1628 -1289
<< locali >>
rect 66 730 118 847
rect 250 730 302 847
rect 150 564 218 598
rect 75 481 218 515
rect 75 315 218 349
rect 150 232 218 266
rect 66 -17 118 100
rect 250 -17 302 100
<< metal1 >>
rect -17 804 385 856
rect 60 306 124 524
rect 152 223 216 607
rect -17 -26 385 26
use nmos130_fast_boundary  MN0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363493
transform 1 0 0 0 1 0
box 0 -84 92 280
use nmos130_fast_boundary  MN0_IBNDR0
timestamp 1704363493
transform 1 0 276 0 1 0
box 0 -84 92 280
use nmos130_fast_center_nf2  MN0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704390143
transform 1 0 92 0 1 0
box -31 -84 215 362
use via_M1_M2_0  MN0_IVD0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704392934
transform 1 0 184 0 1 249
box -17 -17 17 17
use via_M1_M2_0  MN0_IVG0
timestamp 1704392934
transform 1 0 184 0 1 332
box -17 -17 17 17
use via_M1_M2_1  MN0_IVTIED0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 184 0 0 415
timestamp 1704386328
transform 1 0 92 0 1 0
box -26 -26 26 26
use pmos130_fast_boundary  MP0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363574
transform 1 0 0 0 -1 830
box 0 -66 168 369
use pmos130_fast_boundary  MP0_IBNDR0
timestamp 1704363574
transform 1 0 276 0 -1 830
box 0 -66 168 369
use pmos130_fast_center_nf2  MP0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704364343
transform 1 0 92 0 -1 830
box -31 -66 215 369
use via_M1_M2_0  MP0_IVD0
timestamp 1704392934
transform 1 0 184 0 -1 581
box -17 -17 17 17
use via_M1_M2_0  MP0_IVG0
timestamp 1704392934
transform 1 0 184 0 -1 498
box -17 -17 17 17
use via_M1_M2_1  MP0_IVTIED0
array 0 1 184 0 0 -415
timestamp 1704386328
transform 1 0 92 0 -1 830
box -26 -26 26 26
use via_M2_M3_0  NoName_1 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704386899
transform 1 0 92 0 1 332
box -32 -17 32 17
use via_M2_M3_0  NoName_3
timestamp 1704386899
transform 1 0 92 0 1 498
box -32 -17 32 17
use via_M2_M3_0  NoName_5
timestamp 1704386899
transform 1 0 184 0 1 249
box -32 -17 32 17
use via_M2_M3_0  NoName_7
timestamp 1704386899
transform 1 0 184 0 1 581
box -32 -17 32 17
<< labels >>
flabel metal1 92 415 92 415 0 FreeSans 512 90 0 0 I
port 1 nsew
flabel metal1 184 415 184 415 0 FreeSans 512 90 0 0 O
port 2 nsew
flabel metal1 184 830 184 830 0 FreeSans 416 0 0 0 VDD
port 3 nsew
flabel metal1 184 0 184 0 0 FreeSans 416 0 0 0 VSS
port 4 nsew
<< end >>
