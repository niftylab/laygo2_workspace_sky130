magic
tech sky130A
magscale 1 2
timestamp 1679560817
<< checkpaint >>
rect -1300 -1325 6732 3337
<< metal1 >>
rect 114 1688 174 2056
rect 402 1688 462 2056
rect 114 -40 174 328
rect 402 -40 462 328
<< metal2 >>
rect -40 1956 5472 2076
rect 108 1554 468 1614
rect 108 1266 468 1326
rect 108 690 468 750
rect 108 402 468 462
rect -40 -60 5472 60
<< metal3 >>
rect 114 690 174 1326
rect 258 402 318 1614
rect 546 432 606 1584
rect 834 432 894 1584
rect 1122 432 1182 1584
rect 1410 432 1470 1584
rect 1698 432 1758 1584
rect 1986 432 2046 1584
rect 2274 432 2334 1584
rect 2562 432 2622 1584
rect 3426 432 3486 1584
rect 4578 432 4638 1584
rect 5154 432 5214 1584
use nmos13_fast_boundary  MN0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 144 1008
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 432 0 1 0
box 0 0 144 1008
use nmos13_fast_center_nf2  MN0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654175211
transform 1 0 144 0 1 0
box -92 286 380 756
use via_M1_M2_0  MN0_IVD0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 288 0 1 432
box -32 -32 32 32
use via_M1_M2_0  MN0_IVG0
timestamp 1647525606
transform 1 0 288 0 1 720
box -32 -32 32 32
use via_M1_M2_1  MN0_IVTIED0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 288 0 0 1008
timestamp 1647525606
transform 1 0 144 0 1 0
box -32 -32 32 32
use pmos13_fast_boundary  MP0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 2016
box 0 0 144 1008
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 432 0 -1 2016
box 0 0 144 1008
use pmos13_fast_center_nf2  MP0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654091791
transform 1 0 144 0 -1 2016
box -92 132 380 756
use via_M1_M2_0  MP0_IVD0
timestamp 1647525606
transform 1 0 288 0 -1 1584
box -32 -32 32 32
use via_M1_M2_0  MP0_IVG0
timestamp 1647525606
transform 1 0 288 0 -1 1296
box -32 -32 32 32
use via_M1_M2_1  MP0_IVTIED0
array 0 1 288 0 0 -1008
timestamp 1647525606
transform 1 0 144 0 -1 2016
box -32 -32 32 32
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 144 0 1 720
box -38 -38 38 38
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 144 0 1 1296
box -38 -38 38 38
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 288 0 1 432
box -38 -38 38 38
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 288 0 1 1584
box -38 -38 38 38
<< labels >>
flabel metal3 144 1008 144 1008 0 FreeSans 480 90 0 0 I
port 13 nsew
flabel metal3 288 1008 288 1008 0 FreeSans 480 90 0 0 O
port 14 nsew
flabel metal3 576 1008 576 1008 0 FreeSans 480 90 0 0 O
port 15 nsew
flabel metal3 864 1008 864 1008 0 FreeSans 480 90 0 0 O
port 16 nsew
flabel metal3 1152 1008 1152 1008 0 FreeSans 480 90 0 0 O
port 17 nsew
flabel metal3 1440 1008 1440 1008 0 FreeSans 480 90 0 0 O
port 18 nsew
flabel metal3 1728 1008 1728 1008 0 FreeSans 480 90 0 0 O
port 19 nsew
flabel metal3 2016 1008 2016 1008 0 FreeSans 480 90 0 0 O
port 20 nsew
flabel metal3 2304 1008 2304 1008 0 FreeSans 480 90 0 0 O
port 21 nsew
flabel metal3 2592 1008 2592 1008 0 FreeSans 480 90 0 0 O
port 22 nsew
flabel metal3 3456 1008 3456 1008 0 FreeSans 480 90 0 0 O
port 23 nsew
flabel metal3 4608 1008 4608 1008 0 FreeSans 480 90 0 0 O
port 24 nsew
flabel metal3 5184 1008 5184 1008 0 FreeSans 480 90 0 0 O
port 25 nsew
flabel metal3 288 1008 288 1008 0 FreeSans 480 90 0 0 O:
port 26 nsew
flabel metal2 432 2016 432 2016 0 FreeSans 960 0 0 0 VDD
port 28 nsew
flabel metal2 576 2016 576 2016 0 FreeSans 960 0 0 0 VDD
port 29 nsew
flabel metal2 720 2016 720 2016 0 FreeSans 960 0 0 0 VDD
port 30 nsew
flabel metal2 864 2016 864 2016 0 FreeSans 960 0 0 0 VDD
port 31 nsew
flabel metal2 1008 2016 1008 2016 0 FreeSans 960 0 0 0 VDD
port 32 nsew
flabel metal2 1152 2016 1152 2016 0 FreeSans 960 0 0 0 VDD
port 33 nsew
flabel metal2 1296 2016 1296 2016 0 FreeSans 960 0 0 0 VDD
port 34 nsew
flabel metal2 1440 2016 1440 2016 0 FreeSans 960 0 0 0 VDD
port 35 nsew
flabel metal2 1872 2016 1872 2016 0 FreeSans 960 0 0 0 VDD
port 36 nsew
flabel metal2 2448 2016 2448 2016 0 FreeSans 960 0 0 0 VDD
port 37 nsew
flabel metal2 2736 2016 2736 2016 0 FreeSans 960 0 0 0 VDD
port 38 nsew
flabel metal2 288 2016 288 2016 0 FreeSans 960 0 0 0 VDD
port 39 nsew
flabel metal2 432 0 432 0 0 FreeSans 960 0 0 0 VSS
port 41 nsew
flabel metal2 576 0 576 0 0 FreeSans 960 0 0 0 VSS
port 42 nsew
flabel metal2 720 0 720 0 0 FreeSans 960 0 0 0 VSS
port 43 nsew
flabel metal2 864 0 864 0 0 FreeSans 960 0 0 0 VSS
port 44 nsew
flabel metal2 1008 0 1008 0 0 FreeSans 960 0 0 0 VSS
port 45 nsew
flabel metal2 1152 0 1152 0 0 FreeSans 960 0 0 0 VSS
port 46 nsew
flabel metal2 1296 0 1296 0 0 FreeSans 960 0 0 0 VSS
port 47 nsew
flabel metal2 1440 0 1440 0 0 FreeSans 960 0 0 0 VSS
port 48 nsew
flabel metal2 1872 0 1872 0 0 FreeSans 960 0 0 0 VSS
port 49 nsew
flabel metal2 2448 0 2448 0 0 FreeSans 960 0 0 0 VSS
port 50 nsew
flabel metal2 2736 0 2736 0 0 FreeSans 960 0 0 0 VSS
port 51 nsew
flabel metal2 288 0 288 0 0 FreeSans 960 0 0 0 VSS
port 52 nsew
<< end >>
