magic
tech sky130A
timestamp 1679560963
<< checkpaint >>
rect -650 -660 1946 1668
<< metal1 >>
rect 57 844 87 1028
rect 201 844 231 1028
rect 345 844 375 1028
rect 489 844 519 1028
rect 633 844 663 1028
rect 777 844 807 1028
rect 921 844 951 1028
rect 1065 844 1095 1028
rect 1209 844 1239 1028
rect 57 -20 87 164
rect 201 -20 231 164
rect 345 -20 375 164
<< metal2 >>
rect -20 978 1316 1038
rect 106 777 1190 807
rect 106 633 326 663
rect 538 633 758 663
rect 970 633 1190 663
rect 106 345 326 375
rect 538 345 758 375
rect 970 345 1190 375
rect 106 201 830 231
rect 970 201 1190 231
rect 538 129 1262 159
rect -20 -30 1316 30
<< metal3 >>
rect 129 345 159 663
rect 561 345 591 663
rect 993 345 1023 663
rect 1137 201 1167 807
use nmos13_fast_boundary  MN0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 360 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1654175211
transform 1 0 72 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN0_IVD0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 144 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN0_IVG0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 144 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN0_IVTIED0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 2 144 0 0 504
timestamp 1647525606
transform 1 0 72 0 1 0
box -16 -16 16 16
use nmos13_fast_boundary  MN1_IBNDL0
timestamp 1655824928
transform 1 0 432 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN1_IBNDR0
timestamp 1655824928
transform 1 0 792 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN1_IM0
array 0 1 144 0 0 504
timestamp 1654175211
transform 1 0 504 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN1_IVD0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 576 0 1 144
box -16 -16 16 16
use via_M1_M2_0  MN1_IVG0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 576 0 1 360
box -16 -16 16 16
use via_M1_M2_0  MN1_IVS0
array 0 2 144 0 0 504
timestamp 1647525606
transform 1 0 504 0 1 216
box -16 -16 16 16
use nmos13_fast_boundary  MN2_IBNDL0
timestamp 1655824928
transform 1 0 864 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN2_IBNDR0
timestamp 1655824928
transform 1 0 1224 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN2_IM0
array 0 1 144 0 0 504
timestamp 1654175211
transform 1 0 936 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN2_IVD0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 1008 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN2_IVG0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 1008 0 1 360
box -16 -16 16 16
use via_M1_M2_0  MN2_IVS0
array 0 2 144 0 0 504
timestamp 1647525606
transform 1 0 936 0 1 144
box -16 -16 16 16
use pmos13_fast_boundary  MP0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 360 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 -504
timestamp 1654091791
transform 1 0 72 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP0_IVD0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 144 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP0_IVG0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 144 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP0_IVTIED0
array 0 2 144 0 0 -504
timestamp 1647525606
transform 1 0 72 0 -1 1008
box -16 -16 16 16
use pmos13_fast_boundary  MP1_IBNDL0
timestamp 1655825313
transform 1 0 432 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP1_IBNDR0
timestamp 1655825313
transform 1 0 792 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP1_IM0
array 0 1 144 0 0 -504
timestamp 1654091791
transform 1 0 504 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP1_IVD0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 576 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP1_IVG0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 576 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP1_IVTIED0
array 0 2 144 0 0 -504
timestamp 1647525606
transform 1 0 504 0 -1 1008
box -16 -16 16 16
use pmos13_fast_boundary  MP2_IBNDL0
timestamp 1655825313
transform 1 0 864 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP2_IBNDR0
timestamp 1655825313
transform 1 0 1224 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP2_IM0
array 0 1 144 0 0 -504
timestamp 1654091791
transform 1 0 936 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP2_IVD0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 1008 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP2_IVG0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 1008 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP2_IVTIED0
array 0 2 144 0 0 -504
timestamp 1647525606
transform 1 0 936 0 -1 1008
box -16 -16 16 16
use via_M2_M3_0  NoName_0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 1008 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_2
timestamp 1647525786
transform 1 0 1008 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 576 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 576 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_6
timestamp 1647525786
transform 1 0 144 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_8
timestamp 1647525786
transform 1 0 144 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_12
timestamp 1647525786
transform 1 0 1152 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_14
timestamp 1647525786
transform 1 0 1152 0 1 792
box -19 -19 19 19
<< labels >>
flabel metal3 1008 504 1008 504 0 FreeSans 240 90 0 0 A
port 1 nsew
flabel metal3 576 504 576 504 0 FreeSans 240 90 0 0 B
port 2 nsew
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 C
port 3 nsew
flabel metal2 648 1008 648 1008 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel metal2 648 0 648 0 0 FreeSans 480 0 0 0 VSS
port 5 nsew
flabel metal3 1152 504 1152 504 0 FreeSans 240 90 0 0 Y
port 6 nsew
<< end >>
