magic
tech sky130A
magscale 1 2
timestamp 1704363589
<< nwell >>
rect 0 -66 184 369
<< properties >>
string FIXED_BBOX 0 0 184 414
<< end >>
