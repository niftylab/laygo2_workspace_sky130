magic
tech sky130A
timestamp 1679560854
<< checkpaint >>
rect -650 -660 3242 1668
<< metal2 >>
rect -20 978 2612 1038
rect 1137 489 1383 519
rect -20 -30 2612 30
<< metal3 >>
rect 57 360 87 648
rect 1137 201 1167 519
rect 1353 345 1383 519
rect 2433 216 2463 792
use logic_generated_inv_16x  inv0 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 0 0 1 0
box -20 -30 1316 1038
use logic_generated_inv_16x  inv1
timestamp 1679560816
transform 1 0 1296 0 1 0
box -20 -30 1316 1038
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 1152 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 1368 0 1 504
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 I
port 1 nsew
flabel metal3 2448 504 2448 504 0 FreeSans 240 90 0 0 O
port 2 nsew
flabel metal2 1296 1008 1296 1008 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal2 1296 0 1296 0 0 FreeSans 480 0 0 0 VSS
port 4 nsew
<< end >>
