magic
tech sky130A
magscale 1 2
timestamp 1706519206
<< checkpaint >>
rect -1260 -1344 1352 1194
<< pwell >>
rect 0 -84 92 369
<< properties >>
string FIXED_BBOX 0 0 92 414
<< end >>
