magic
tech sky130A
timestamp 1655825501
<< nwell >>
rect 0 66 72 342
<< labels >>
flabel space 0 0 72 512 0 FreeSans 160 90 0 0 PTAP_LEFT
<< end >>
