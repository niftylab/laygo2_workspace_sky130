magic
tech sky130A
timestamp 1655825515
<< checkpaint >>
rect -630 -526 702 854
<< nwell >>
rect 0 66 72 342
<< labels >>
flabel space 0 0 72 315 0 FreeSans 160 90 0 0 PTAP_RIGHT
<< end >>
