magic
tech sky130A
magscale 1 2
timestamp 1668535077
<< nwell >>
rect 0 3348 21024 3900
rect 0 132 21024 684
<< pwell >>
rect 0 2388 21024 2700
rect 0 1332 21024 1644
<< pmos >>
rect 778 3384 808 3864
rect 922 3384 952 3864
rect 1354 3384 1384 3864
rect 1498 3384 1528 3864
rect 1930 3384 1960 3864
rect 2074 3384 2104 3864
rect 2506 3384 2536 3864
rect 2650 3384 2680 3864
rect 3080 3384 3110 3864
rect 3224 3384 3254 3864
rect 4232 3384 4262 3864
rect 4376 3384 4406 3864
rect 4808 3384 4838 3864
rect 4952 3384 4982 3864
rect 5384 3384 5414 3864
rect 5528 3384 5558 3864
rect 5960 3384 5990 3864
rect 6104 3384 6134 3864
rect 6536 3384 6566 3864
rect 6680 3384 6710 3864
rect 7688 3384 7718 3864
rect 7832 3384 7862 3864
rect 8264 3384 8294 3864
rect 8408 3384 8438 3864
rect 8840 3384 8870 3864
rect 8984 3384 9014 3864
rect 9416 3384 9446 3864
rect 9560 3384 9590 3864
rect 10280 3384 10310 3864
rect 10424 3384 10454 3864
rect 10856 3384 10886 3864
rect 11000 3384 11030 3864
rect 12008 3384 12038 3864
rect 12152 3384 12182 3864
rect 12584 3384 12614 3864
rect 12728 3384 12758 3864
rect 13736 3384 13766 3864
rect 13880 3384 13910 3864
rect 14312 3384 14342 3864
rect 14456 3384 14486 3864
rect 14888 3384 14918 3864
rect 15032 3384 15062 3864
rect 16618 3384 16648 3864
rect 16762 3384 16792 3864
rect 16906 3384 16936 3864
rect 17050 3384 17080 3864
rect 17194 3384 17224 3864
rect 17338 3384 17368 3864
rect 17482 3384 17512 3864
rect 17626 3384 17656 3864
rect 17770 3384 17800 3864
rect 17914 3384 17944 3864
rect 18058 3384 18088 3864
rect 18202 3384 18232 3864
rect 18346 3384 18376 3864
rect 18490 3384 18520 3864
rect 18634 3384 18664 3864
rect 18778 3384 18808 3864
rect 18922 3384 18952 3864
rect 19066 3384 19096 3864
rect 19210 3384 19240 3864
rect 19354 3384 19384 3864
rect 19498 3384 19528 3864
rect 19642 3384 19672 3864
rect 19786 3384 19816 3864
rect 19930 3384 19960 3864
rect 776 168 806 648
rect 920 168 950 648
rect 1352 168 1382 648
rect 1496 168 1526 648
rect 1928 168 1958 648
rect 2072 168 2102 648
rect 3080 168 3110 648
rect 3224 168 3254 648
rect 3656 168 3686 648
rect 3800 168 3830 648
rect 4232 168 4262 648
rect 4376 168 4406 648
rect 5960 168 5990 648
rect 6104 168 6134 648
rect 6536 168 6566 648
rect 6680 168 6710 648
rect 7112 168 7142 648
rect 7256 168 7286 648
rect 7688 168 7718 648
rect 7832 168 7862 648
rect 8264 168 8294 648
rect 8408 168 8438 648
rect 9416 168 9446 648
rect 9560 168 9590 648
rect 9992 168 10022 648
rect 10136 168 10166 648
rect 10568 168 10598 648
rect 10712 168 10742 648
rect 11144 168 11174 648
rect 11288 168 11318 648
rect 12008 168 12038 648
rect 12152 168 12182 648
rect 12584 168 12614 648
rect 12728 168 12758 648
rect 13160 168 13190 648
rect 13304 168 13334 648
rect 13736 168 13766 648
rect 13880 168 13910 648
rect 14888 168 14918 648
rect 15032 168 15062 648
rect 15466 168 15496 648
rect 15610 168 15640 648
rect 16040 168 16070 648
rect 16184 168 16214 648
rect 16328 168 16358 648
rect 16472 168 16502 648
rect 17480 168 17510 648
rect 17624 168 17654 648
rect 17768 168 17798 648
rect 17912 168 17942 648
rect 18056 168 18086 648
rect 18200 168 18230 648
rect 18344 168 18374 648
rect 18488 168 18518 648
rect 18632 168 18662 648
rect 18776 168 18806 648
rect 18920 168 18950 648
rect 19064 168 19094 648
rect 19208 168 19238 648
rect 19352 168 19382 648
rect 19496 168 19526 648
rect 19640 168 19670 648
rect 19784 168 19814 648
rect 19928 168 19958 648
rect 20072 168 20102 648
rect 20216 168 20246 648
rect 20360 168 20390 648
rect 20504 168 20534 648
rect 20648 168 20678 648
rect 20792 168 20822 648
<< nmoslvt >>
rect 778 2424 808 2664
rect 922 2424 952 2664
rect 1354 2424 1384 2664
rect 1498 2424 1528 2664
rect 1930 2424 1960 2664
rect 2074 2424 2104 2664
rect 2506 2424 2536 2664
rect 2650 2424 2680 2664
rect 3080 2424 3110 2664
rect 3224 2424 3254 2664
rect 4232 2424 4262 2664
rect 4376 2424 4406 2664
rect 4808 2424 4838 2664
rect 4952 2424 4982 2664
rect 5384 2424 5414 2664
rect 5528 2424 5558 2664
rect 5960 2424 5990 2664
rect 6104 2424 6134 2664
rect 6536 2424 6566 2664
rect 6680 2424 6710 2664
rect 7688 2424 7718 2664
rect 7832 2424 7862 2664
rect 8264 2424 8294 2664
rect 8408 2424 8438 2664
rect 8840 2424 8870 2664
rect 8984 2424 9014 2664
rect 9416 2424 9446 2664
rect 9560 2424 9590 2664
rect 10280 2424 10310 2664
rect 10424 2424 10454 2664
rect 10856 2424 10886 2664
rect 11000 2424 11030 2664
rect 12008 2424 12038 2664
rect 12152 2424 12182 2664
rect 12584 2424 12614 2664
rect 12728 2424 12758 2664
rect 13736 2424 13766 2664
rect 13880 2424 13910 2664
rect 14312 2424 14342 2664
rect 14456 2424 14486 2664
rect 14888 2424 14918 2664
rect 15032 2424 15062 2664
rect 16618 2424 16648 2664
rect 16762 2424 16792 2664
rect 16906 2424 16936 2664
rect 17050 2424 17080 2664
rect 17194 2424 17224 2664
rect 17338 2424 17368 2664
rect 17482 2424 17512 2664
rect 17626 2424 17656 2664
rect 17770 2424 17800 2664
rect 17914 2424 17944 2664
rect 18058 2424 18088 2664
rect 18202 2424 18232 2664
rect 18346 2424 18376 2664
rect 18490 2424 18520 2664
rect 18634 2424 18664 2664
rect 18778 2424 18808 2664
rect 18922 2424 18952 2664
rect 19066 2424 19096 2664
rect 19210 2424 19240 2664
rect 19354 2424 19384 2664
rect 19498 2424 19528 2664
rect 19642 2424 19672 2664
rect 19786 2424 19816 2664
rect 19930 2424 19960 2664
rect 776 1368 806 1608
rect 920 1368 950 1608
rect 1352 1368 1382 1608
rect 1496 1368 1526 1608
rect 1928 1368 1958 1608
rect 2072 1368 2102 1608
rect 3080 1368 3110 1608
rect 3224 1368 3254 1608
rect 3656 1368 3686 1608
rect 3800 1368 3830 1608
rect 4232 1368 4262 1608
rect 4376 1368 4406 1608
rect 5960 1368 5990 1608
rect 6104 1368 6134 1608
rect 6536 1368 6566 1608
rect 6680 1368 6710 1608
rect 7112 1368 7142 1608
rect 7256 1368 7286 1608
rect 7688 1368 7718 1608
rect 7832 1368 7862 1608
rect 8264 1368 8294 1608
rect 8408 1368 8438 1608
rect 9416 1368 9446 1608
rect 9560 1368 9590 1608
rect 9992 1368 10022 1608
rect 10136 1368 10166 1608
rect 10568 1368 10598 1608
rect 10712 1368 10742 1608
rect 11144 1368 11174 1608
rect 11288 1368 11318 1608
rect 12008 1368 12038 1608
rect 12152 1368 12182 1608
rect 12584 1368 12614 1608
rect 12728 1368 12758 1608
rect 13160 1368 13190 1608
rect 13304 1368 13334 1608
rect 13736 1368 13766 1608
rect 13880 1368 13910 1608
rect 14888 1368 14918 1608
rect 15032 1368 15062 1608
rect 15466 1368 15496 1608
rect 15610 1368 15640 1608
rect 16040 1368 16070 1608
rect 16184 1368 16214 1608
rect 16328 1368 16358 1608
rect 16472 1368 16502 1608
rect 17480 1368 17510 1608
rect 17624 1368 17654 1608
rect 17768 1368 17798 1608
rect 17912 1368 17942 1608
rect 18056 1368 18086 1608
rect 18200 1368 18230 1608
rect 18344 1368 18374 1608
rect 18488 1368 18518 1608
rect 18632 1368 18662 1608
rect 18776 1368 18806 1608
rect 18920 1368 18950 1608
rect 19064 1368 19094 1608
rect 19208 1368 19238 1608
rect 19352 1368 19382 1608
rect 19496 1368 19526 1608
rect 19640 1368 19670 1608
rect 19784 1368 19814 1608
rect 19928 1368 19958 1608
rect 20072 1368 20102 1608
rect 20216 1368 20246 1608
rect 20360 1368 20390 1608
rect 20504 1368 20534 1608
rect 20648 1368 20678 1608
rect 20792 1368 20822 1608
<< ndiff >>
rect 664 2614 778 2664
rect 664 2574 700 2614
rect 740 2574 778 2614
rect 664 2514 778 2574
rect 664 2474 700 2514
rect 740 2474 778 2514
rect 664 2424 778 2474
rect 808 2614 922 2664
rect 808 2574 844 2614
rect 884 2574 922 2614
rect 808 2514 922 2574
rect 808 2474 844 2514
rect 884 2474 922 2514
rect 808 2424 922 2474
rect 952 2614 1064 2664
rect 952 2574 988 2614
rect 1028 2574 1064 2614
rect 952 2514 1064 2574
rect 952 2474 988 2514
rect 1028 2474 1064 2514
rect 952 2424 1064 2474
rect 1240 2614 1354 2664
rect 1240 2574 1276 2614
rect 1316 2574 1354 2614
rect 1240 2514 1354 2574
rect 1240 2474 1276 2514
rect 1316 2474 1354 2514
rect 1240 2424 1354 2474
rect 1384 2614 1498 2664
rect 1384 2574 1420 2614
rect 1460 2574 1498 2614
rect 1384 2514 1498 2574
rect 1384 2474 1420 2514
rect 1460 2474 1498 2514
rect 1384 2424 1498 2474
rect 1528 2614 1640 2664
rect 1528 2574 1564 2614
rect 1604 2574 1640 2614
rect 1528 2514 1640 2574
rect 1528 2474 1564 2514
rect 1604 2474 1640 2514
rect 1528 2424 1640 2474
rect 1816 2614 1930 2664
rect 1816 2574 1852 2614
rect 1892 2574 1930 2614
rect 1816 2514 1930 2574
rect 1816 2474 1852 2514
rect 1892 2474 1930 2514
rect 1816 2424 1930 2474
rect 1960 2614 2074 2664
rect 1960 2574 1996 2614
rect 2036 2574 2074 2614
rect 1960 2514 2074 2574
rect 1960 2474 1996 2514
rect 2036 2474 2074 2514
rect 1960 2424 2074 2474
rect 2104 2614 2216 2664
rect 2104 2574 2140 2614
rect 2180 2574 2216 2614
rect 2104 2514 2216 2574
rect 2104 2474 2140 2514
rect 2180 2474 2216 2514
rect 2104 2424 2216 2474
rect 2392 2614 2506 2664
rect 2392 2574 2428 2614
rect 2468 2574 2506 2614
rect 2392 2514 2506 2574
rect 2392 2474 2428 2514
rect 2468 2474 2506 2514
rect 2392 2424 2506 2474
rect 2536 2614 2650 2664
rect 2536 2574 2572 2614
rect 2612 2574 2650 2614
rect 2536 2514 2650 2574
rect 2536 2474 2572 2514
rect 2612 2474 2650 2514
rect 2536 2424 2650 2474
rect 2680 2614 2792 2664
rect 2680 2574 2716 2614
rect 2756 2574 2792 2614
rect 2680 2514 2792 2574
rect 2680 2474 2716 2514
rect 2756 2474 2792 2514
rect 2680 2424 2792 2474
rect 2968 2614 3080 2664
rect 2968 2574 3004 2614
rect 3044 2574 3080 2614
rect 2968 2514 3080 2574
rect 2968 2474 3004 2514
rect 3044 2474 3080 2514
rect 2968 2424 3080 2474
rect 3110 2614 3224 2664
rect 3110 2574 3148 2614
rect 3188 2574 3224 2614
rect 3110 2514 3224 2574
rect 3110 2474 3148 2514
rect 3188 2474 3224 2514
rect 3110 2424 3224 2474
rect 3254 2614 3368 2664
rect 3254 2574 3292 2614
rect 3332 2574 3368 2614
rect 3254 2514 3368 2574
rect 3254 2474 3292 2514
rect 3332 2474 3368 2514
rect 3254 2424 3368 2474
rect 4120 2614 4232 2664
rect 4120 2574 4156 2614
rect 4196 2574 4232 2614
rect 4120 2514 4232 2574
rect 4120 2474 4156 2514
rect 4196 2474 4232 2514
rect 4120 2424 4232 2474
rect 4262 2614 4376 2664
rect 4262 2574 4300 2614
rect 4340 2574 4376 2614
rect 4262 2514 4376 2574
rect 4262 2474 4300 2514
rect 4340 2474 4376 2514
rect 4262 2424 4376 2474
rect 4406 2614 4520 2664
rect 4406 2574 4444 2614
rect 4484 2574 4520 2614
rect 4406 2514 4520 2574
rect 4406 2474 4444 2514
rect 4484 2474 4520 2514
rect 4406 2424 4520 2474
rect 4696 2614 4808 2664
rect 4696 2574 4732 2614
rect 4772 2574 4808 2614
rect 4696 2514 4808 2574
rect 4696 2474 4732 2514
rect 4772 2474 4808 2514
rect 4696 2424 4808 2474
rect 4838 2614 4952 2664
rect 4838 2574 4876 2614
rect 4916 2574 4952 2614
rect 4838 2514 4952 2574
rect 4838 2474 4876 2514
rect 4916 2474 4952 2514
rect 4838 2424 4952 2474
rect 4982 2614 5096 2664
rect 4982 2574 5020 2614
rect 5060 2574 5096 2614
rect 4982 2514 5096 2574
rect 4982 2474 5020 2514
rect 5060 2474 5096 2514
rect 4982 2424 5096 2474
rect 5272 2614 5384 2664
rect 5272 2574 5308 2614
rect 5348 2574 5384 2614
rect 5272 2514 5384 2574
rect 5272 2474 5308 2514
rect 5348 2474 5384 2514
rect 5272 2424 5384 2474
rect 5414 2614 5528 2664
rect 5414 2574 5452 2614
rect 5492 2574 5528 2614
rect 5414 2514 5528 2574
rect 5414 2474 5452 2514
rect 5492 2474 5528 2514
rect 5414 2424 5528 2474
rect 5558 2614 5672 2664
rect 5558 2574 5596 2614
rect 5636 2574 5672 2614
rect 5558 2514 5672 2574
rect 5558 2474 5596 2514
rect 5636 2474 5672 2514
rect 5558 2424 5672 2474
rect 5848 2614 5960 2664
rect 5848 2574 5884 2614
rect 5924 2574 5960 2614
rect 5848 2514 5960 2574
rect 5848 2474 5884 2514
rect 5924 2474 5960 2514
rect 5848 2424 5960 2474
rect 5990 2614 6104 2664
rect 5990 2574 6028 2614
rect 6068 2574 6104 2614
rect 5990 2514 6104 2574
rect 5990 2474 6028 2514
rect 6068 2474 6104 2514
rect 5990 2424 6104 2474
rect 6134 2614 6248 2664
rect 6134 2574 6172 2614
rect 6212 2574 6248 2614
rect 6134 2514 6248 2574
rect 6134 2474 6172 2514
rect 6212 2474 6248 2514
rect 6134 2424 6248 2474
rect 6424 2614 6536 2664
rect 6424 2574 6460 2614
rect 6500 2574 6536 2614
rect 6424 2514 6536 2574
rect 6424 2474 6460 2514
rect 6500 2474 6536 2514
rect 6424 2424 6536 2474
rect 6566 2614 6680 2664
rect 6566 2574 6604 2614
rect 6644 2574 6680 2614
rect 6566 2514 6680 2574
rect 6566 2474 6604 2514
rect 6644 2474 6680 2514
rect 6566 2424 6680 2474
rect 6710 2614 6824 2664
rect 6710 2574 6748 2614
rect 6788 2574 6824 2614
rect 6710 2514 6824 2574
rect 6710 2474 6748 2514
rect 6788 2474 6824 2514
rect 6710 2424 6824 2474
rect 7576 2614 7688 2664
rect 7576 2574 7612 2614
rect 7652 2574 7688 2614
rect 7576 2514 7688 2574
rect 7576 2474 7612 2514
rect 7652 2474 7688 2514
rect 7576 2424 7688 2474
rect 7718 2614 7832 2664
rect 7718 2574 7756 2614
rect 7796 2574 7832 2614
rect 7718 2514 7832 2574
rect 7718 2474 7756 2514
rect 7796 2474 7832 2514
rect 7718 2424 7832 2474
rect 7862 2614 7976 2664
rect 7862 2574 7900 2614
rect 7940 2574 7976 2614
rect 7862 2514 7976 2574
rect 7862 2474 7900 2514
rect 7940 2474 7976 2514
rect 7862 2424 7976 2474
rect 8152 2614 8264 2664
rect 8152 2574 8188 2614
rect 8228 2574 8264 2614
rect 8152 2514 8264 2574
rect 8152 2474 8188 2514
rect 8228 2474 8264 2514
rect 8152 2424 8264 2474
rect 8294 2614 8408 2664
rect 8294 2574 8332 2614
rect 8372 2574 8408 2614
rect 8294 2514 8408 2574
rect 8294 2474 8332 2514
rect 8372 2474 8408 2514
rect 8294 2424 8408 2474
rect 8438 2614 8552 2664
rect 8438 2574 8476 2614
rect 8516 2574 8552 2614
rect 8438 2514 8552 2574
rect 8438 2474 8476 2514
rect 8516 2474 8552 2514
rect 8438 2424 8552 2474
rect 8728 2614 8840 2664
rect 8728 2574 8764 2614
rect 8804 2574 8840 2614
rect 8728 2514 8840 2574
rect 8728 2474 8764 2514
rect 8804 2474 8840 2514
rect 8728 2424 8840 2474
rect 8870 2614 8984 2664
rect 8870 2574 8908 2614
rect 8948 2574 8984 2614
rect 8870 2514 8984 2574
rect 8870 2474 8908 2514
rect 8948 2474 8984 2514
rect 8870 2424 8984 2474
rect 9014 2614 9128 2664
rect 9014 2574 9052 2614
rect 9092 2574 9128 2614
rect 9014 2514 9128 2574
rect 9014 2474 9052 2514
rect 9092 2474 9128 2514
rect 9014 2424 9128 2474
rect 9304 2614 9416 2664
rect 9304 2574 9340 2614
rect 9380 2574 9416 2614
rect 9304 2514 9416 2574
rect 9304 2474 9340 2514
rect 9380 2474 9416 2514
rect 9304 2424 9416 2474
rect 9446 2614 9560 2664
rect 9446 2574 9484 2614
rect 9524 2574 9560 2614
rect 9446 2514 9560 2574
rect 9446 2474 9484 2514
rect 9524 2474 9560 2514
rect 9446 2424 9560 2474
rect 9590 2614 9704 2664
rect 9590 2574 9628 2614
rect 9668 2574 9704 2614
rect 9590 2514 9704 2574
rect 9590 2474 9628 2514
rect 9668 2474 9704 2514
rect 9590 2424 9704 2474
rect 10168 2614 10280 2664
rect 10168 2574 10204 2614
rect 10244 2574 10280 2614
rect 10168 2514 10280 2574
rect 10168 2474 10204 2514
rect 10244 2474 10280 2514
rect 10168 2424 10280 2474
rect 10310 2614 10424 2664
rect 10310 2574 10348 2614
rect 10388 2574 10424 2614
rect 10310 2514 10424 2574
rect 10310 2474 10348 2514
rect 10388 2474 10424 2514
rect 10310 2424 10424 2474
rect 10454 2614 10568 2664
rect 10454 2574 10492 2614
rect 10532 2574 10568 2614
rect 10454 2514 10568 2574
rect 10454 2474 10492 2514
rect 10532 2474 10568 2514
rect 10454 2424 10568 2474
rect 10744 2614 10856 2664
rect 10744 2574 10780 2614
rect 10820 2574 10856 2614
rect 10744 2514 10856 2574
rect 10744 2474 10780 2514
rect 10820 2474 10856 2514
rect 10744 2424 10856 2474
rect 10886 2614 11000 2664
rect 10886 2574 10924 2614
rect 10964 2574 11000 2614
rect 10886 2514 11000 2574
rect 10886 2474 10924 2514
rect 10964 2474 11000 2514
rect 10886 2424 11000 2474
rect 11030 2614 11144 2664
rect 11030 2574 11068 2614
rect 11108 2574 11144 2614
rect 11030 2514 11144 2574
rect 11030 2474 11068 2514
rect 11108 2474 11144 2514
rect 11030 2424 11144 2474
rect 11896 2614 12008 2664
rect 11896 2574 11932 2614
rect 11972 2574 12008 2614
rect 11896 2514 12008 2574
rect 11896 2474 11932 2514
rect 11972 2474 12008 2514
rect 11896 2424 12008 2474
rect 12038 2614 12152 2664
rect 12038 2574 12076 2614
rect 12116 2574 12152 2614
rect 12038 2514 12152 2574
rect 12038 2474 12076 2514
rect 12116 2474 12152 2514
rect 12038 2424 12152 2474
rect 12182 2614 12296 2664
rect 12182 2574 12220 2614
rect 12260 2574 12296 2614
rect 12182 2514 12296 2574
rect 12182 2474 12220 2514
rect 12260 2474 12296 2514
rect 12182 2424 12296 2474
rect 12472 2614 12584 2664
rect 12472 2574 12508 2614
rect 12548 2574 12584 2614
rect 12472 2514 12584 2574
rect 12472 2474 12508 2514
rect 12548 2474 12584 2514
rect 12472 2424 12584 2474
rect 12614 2614 12728 2664
rect 12614 2574 12652 2614
rect 12692 2574 12728 2614
rect 12614 2514 12728 2574
rect 12614 2474 12652 2514
rect 12692 2474 12728 2514
rect 12614 2424 12728 2474
rect 12758 2614 12872 2664
rect 12758 2574 12796 2614
rect 12836 2574 12872 2614
rect 12758 2514 12872 2574
rect 12758 2474 12796 2514
rect 12836 2474 12872 2514
rect 12758 2424 12872 2474
rect 13624 2614 13736 2664
rect 13624 2574 13660 2614
rect 13700 2574 13736 2614
rect 13624 2514 13736 2574
rect 13624 2474 13660 2514
rect 13700 2474 13736 2514
rect 13624 2424 13736 2474
rect 13766 2614 13880 2664
rect 13766 2574 13804 2614
rect 13844 2574 13880 2614
rect 13766 2514 13880 2574
rect 13766 2474 13804 2514
rect 13844 2474 13880 2514
rect 13766 2424 13880 2474
rect 13910 2614 14024 2664
rect 13910 2574 13948 2614
rect 13988 2574 14024 2614
rect 13910 2514 14024 2574
rect 13910 2474 13948 2514
rect 13988 2474 14024 2514
rect 13910 2424 14024 2474
rect 14200 2614 14312 2664
rect 14200 2574 14236 2614
rect 14276 2574 14312 2614
rect 14200 2514 14312 2574
rect 14200 2474 14236 2514
rect 14276 2474 14312 2514
rect 14200 2424 14312 2474
rect 14342 2614 14456 2664
rect 14342 2574 14380 2614
rect 14420 2574 14456 2614
rect 14342 2514 14456 2574
rect 14342 2474 14380 2514
rect 14420 2474 14456 2514
rect 14342 2424 14456 2474
rect 14486 2614 14600 2664
rect 14486 2574 14524 2614
rect 14564 2574 14600 2614
rect 14486 2514 14600 2574
rect 14486 2474 14524 2514
rect 14564 2474 14600 2514
rect 14486 2424 14600 2474
rect 14776 2614 14888 2664
rect 14776 2574 14812 2614
rect 14852 2574 14888 2614
rect 14776 2514 14888 2574
rect 14776 2474 14812 2514
rect 14852 2474 14888 2514
rect 14776 2424 14888 2474
rect 14918 2614 15032 2664
rect 14918 2574 14956 2614
rect 14996 2574 15032 2614
rect 14918 2514 15032 2574
rect 14918 2474 14956 2514
rect 14996 2474 15032 2514
rect 14918 2424 15032 2474
rect 15062 2614 15176 2664
rect 15062 2574 15100 2614
rect 15140 2574 15176 2614
rect 15062 2514 15176 2574
rect 15062 2474 15100 2514
rect 15140 2474 15176 2514
rect 15062 2424 15176 2474
rect 16504 2614 16618 2664
rect 16504 2574 16540 2614
rect 16580 2574 16618 2614
rect 16504 2514 16618 2574
rect 16504 2474 16540 2514
rect 16580 2474 16618 2514
rect 16504 2424 16618 2474
rect 16648 2614 16762 2664
rect 16648 2574 16684 2614
rect 16724 2574 16762 2614
rect 16648 2514 16762 2574
rect 16648 2474 16684 2514
rect 16724 2474 16762 2514
rect 16648 2424 16762 2474
rect 16792 2614 16906 2664
rect 16792 2574 16828 2614
rect 16868 2574 16906 2614
rect 16792 2514 16906 2574
rect 16792 2474 16828 2514
rect 16868 2474 16906 2514
rect 16792 2424 16906 2474
rect 16936 2614 17050 2664
rect 16936 2574 16972 2614
rect 17012 2574 17050 2614
rect 16936 2514 17050 2574
rect 16936 2474 16972 2514
rect 17012 2474 17050 2514
rect 16936 2424 17050 2474
rect 17080 2614 17194 2664
rect 17080 2574 17116 2614
rect 17156 2574 17194 2614
rect 17080 2514 17194 2574
rect 17080 2474 17116 2514
rect 17156 2474 17194 2514
rect 17080 2424 17194 2474
rect 17224 2614 17338 2664
rect 17224 2574 17260 2614
rect 17300 2574 17338 2614
rect 17224 2514 17338 2574
rect 17224 2474 17260 2514
rect 17300 2474 17338 2514
rect 17224 2424 17338 2474
rect 17368 2614 17482 2664
rect 17368 2574 17404 2614
rect 17444 2574 17482 2614
rect 17368 2514 17482 2574
rect 17368 2474 17404 2514
rect 17444 2474 17482 2514
rect 17368 2424 17482 2474
rect 17512 2614 17626 2664
rect 17512 2574 17548 2614
rect 17588 2574 17626 2614
rect 17512 2514 17626 2574
rect 17512 2474 17548 2514
rect 17588 2474 17626 2514
rect 17512 2424 17626 2474
rect 17656 2614 17770 2664
rect 17656 2574 17692 2614
rect 17732 2574 17770 2614
rect 17656 2514 17770 2574
rect 17656 2474 17692 2514
rect 17732 2474 17770 2514
rect 17656 2424 17770 2474
rect 17800 2614 17914 2664
rect 17800 2574 17836 2614
rect 17876 2574 17914 2614
rect 17800 2514 17914 2574
rect 17800 2474 17836 2514
rect 17876 2474 17914 2514
rect 17800 2424 17914 2474
rect 17944 2614 18058 2664
rect 17944 2574 17980 2614
rect 18020 2574 18058 2614
rect 17944 2514 18058 2574
rect 17944 2474 17980 2514
rect 18020 2474 18058 2514
rect 17944 2424 18058 2474
rect 18088 2614 18202 2664
rect 18088 2574 18124 2614
rect 18164 2574 18202 2614
rect 18088 2514 18202 2574
rect 18088 2474 18124 2514
rect 18164 2474 18202 2514
rect 18088 2424 18202 2474
rect 18232 2614 18346 2664
rect 18232 2574 18268 2614
rect 18308 2574 18346 2614
rect 18232 2514 18346 2574
rect 18232 2474 18268 2514
rect 18308 2474 18346 2514
rect 18232 2424 18346 2474
rect 18376 2614 18490 2664
rect 18376 2574 18412 2614
rect 18452 2574 18490 2614
rect 18376 2514 18490 2574
rect 18376 2474 18412 2514
rect 18452 2474 18490 2514
rect 18376 2424 18490 2474
rect 18520 2614 18634 2664
rect 18520 2574 18556 2614
rect 18596 2574 18634 2614
rect 18520 2514 18634 2574
rect 18520 2474 18556 2514
rect 18596 2474 18634 2514
rect 18520 2424 18634 2474
rect 18664 2614 18778 2664
rect 18664 2574 18700 2614
rect 18740 2574 18778 2614
rect 18664 2514 18778 2574
rect 18664 2474 18700 2514
rect 18740 2474 18778 2514
rect 18664 2424 18778 2474
rect 18808 2614 18922 2664
rect 18808 2574 18844 2614
rect 18884 2574 18922 2614
rect 18808 2514 18922 2574
rect 18808 2474 18844 2514
rect 18884 2474 18922 2514
rect 18808 2424 18922 2474
rect 18952 2614 19066 2664
rect 18952 2574 18988 2614
rect 19028 2574 19066 2614
rect 18952 2514 19066 2574
rect 18952 2474 18988 2514
rect 19028 2474 19066 2514
rect 18952 2424 19066 2474
rect 19096 2614 19210 2664
rect 19096 2574 19132 2614
rect 19172 2574 19210 2614
rect 19096 2514 19210 2574
rect 19096 2474 19132 2514
rect 19172 2474 19210 2514
rect 19096 2424 19210 2474
rect 19240 2614 19354 2664
rect 19240 2574 19276 2614
rect 19316 2574 19354 2614
rect 19240 2514 19354 2574
rect 19240 2474 19276 2514
rect 19316 2474 19354 2514
rect 19240 2424 19354 2474
rect 19384 2614 19498 2664
rect 19384 2574 19420 2614
rect 19460 2574 19498 2614
rect 19384 2514 19498 2574
rect 19384 2474 19420 2514
rect 19460 2474 19498 2514
rect 19384 2424 19498 2474
rect 19528 2614 19642 2664
rect 19528 2574 19564 2614
rect 19604 2574 19642 2614
rect 19528 2514 19642 2574
rect 19528 2474 19564 2514
rect 19604 2474 19642 2514
rect 19528 2424 19642 2474
rect 19672 2614 19786 2664
rect 19672 2574 19708 2614
rect 19748 2574 19786 2614
rect 19672 2514 19786 2574
rect 19672 2474 19708 2514
rect 19748 2474 19786 2514
rect 19672 2424 19786 2474
rect 19816 2614 19930 2664
rect 19816 2574 19852 2614
rect 19892 2574 19930 2614
rect 19816 2514 19930 2574
rect 19816 2474 19852 2514
rect 19892 2474 19930 2514
rect 19816 2424 19930 2474
rect 19960 2614 20072 2664
rect 19960 2574 19996 2614
rect 20036 2574 20072 2614
rect 19960 2514 20072 2574
rect 19960 2474 19996 2514
rect 20036 2474 20072 2514
rect 19960 2424 20072 2474
rect 664 1558 776 1608
rect 664 1518 700 1558
rect 740 1518 776 1558
rect 664 1458 776 1518
rect 664 1418 700 1458
rect 740 1418 776 1458
rect 664 1368 776 1418
rect 806 1558 920 1608
rect 806 1518 844 1558
rect 884 1518 920 1558
rect 806 1458 920 1518
rect 806 1418 844 1458
rect 884 1418 920 1458
rect 806 1368 920 1418
rect 950 1558 1064 1608
rect 950 1518 988 1558
rect 1028 1518 1064 1558
rect 950 1458 1064 1518
rect 950 1418 988 1458
rect 1028 1418 1064 1458
rect 950 1368 1064 1418
rect 1240 1558 1352 1608
rect 1240 1518 1276 1558
rect 1316 1518 1352 1558
rect 1240 1458 1352 1518
rect 1240 1418 1276 1458
rect 1316 1418 1352 1458
rect 1240 1368 1352 1418
rect 1382 1558 1496 1608
rect 1382 1518 1420 1558
rect 1460 1518 1496 1558
rect 1382 1458 1496 1518
rect 1382 1418 1420 1458
rect 1460 1418 1496 1458
rect 1382 1368 1496 1418
rect 1526 1558 1640 1608
rect 1526 1518 1564 1558
rect 1604 1518 1640 1558
rect 1526 1458 1640 1518
rect 1526 1418 1564 1458
rect 1604 1418 1640 1458
rect 1526 1368 1640 1418
rect 1816 1558 1928 1608
rect 1816 1518 1852 1558
rect 1892 1518 1928 1558
rect 1816 1458 1928 1518
rect 1816 1418 1852 1458
rect 1892 1418 1928 1458
rect 1816 1368 1928 1418
rect 1958 1558 2072 1608
rect 1958 1518 1996 1558
rect 2036 1518 2072 1558
rect 1958 1458 2072 1518
rect 1958 1418 1996 1458
rect 2036 1418 2072 1458
rect 1958 1368 2072 1418
rect 2102 1558 2216 1608
rect 2102 1518 2140 1558
rect 2180 1518 2216 1558
rect 2102 1458 2216 1518
rect 2102 1418 2140 1458
rect 2180 1418 2216 1458
rect 2102 1368 2216 1418
rect 2968 1558 3080 1608
rect 2968 1518 3004 1558
rect 3044 1518 3080 1558
rect 2968 1458 3080 1518
rect 2968 1418 3004 1458
rect 3044 1418 3080 1458
rect 2968 1368 3080 1418
rect 3110 1558 3224 1608
rect 3110 1518 3148 1558
rect 3188 1518 3224 1558
rect 3110 1458 3224 1518
rect 3110 1418 3148 1458
rect 3188 1418 3224 1458
rect 3110 1368 3224 1418
rect 3254 1558 3368 1608
rect 3254 1518 3292 1558
rect 3332 1518 3368 1558
rect 3254 1458 3368 1518
rect 3254 1418 3292 1458
rect 3332 1418 3368 1458
rect 3254 1368 3368 1418
rect 3544 1558 3656 1608
rect 3544 1518 3580 1558
rect 3620 1518 3656 1558
rect 3544 1458 3656 1518
rect 3544 1418 3580 1458
rect 3620 1418 3656 1458
rect 3544 1368 3656 1418
rect 3686 1558 3800 1608
rect 3686 1518 3724 1558
rect 3764 1518 3800 1558
rect 3686 1458 3800 1518
rect 3686 1418 3724 1458
rect 3764 1418 3800 1458
rect 3686 1368 3800 1418
rect 3830 1558 3944 1608
rect 3830 1518 3868 1558
rect 3908 1518 3944 1558
rect 3830 1458 3944 1518
rect 3830 1418 3868 1458
rect 3908 1418 3944 1458
rect 3830 1368 3944 1418
rect 4120 1558 4232 1608
rect 4120 1518 4156 1558
rect 4196 1518 4232 1558
rect 4120 1458 4232 1518
rect 4120 1418 4156 1458
rect 4196 1418 4232 1458
rect 4120 1368 4232 1418
rect 4262 1558 4376 1608
rect 4262 1518 4300 1558
rect 4340 1518 4376 1558
rect 4262 1458 4376 1518
rect 4262 1418 4300 1458
rect 4340 1418 4376 1458
rect 4262 1368 4376 1418
rect 4406 1558 4520 1608
rect 4406 1518 4444 1558
rect 4484 1518 4520 1558
rect 4406 1458 4520 1518
rect 4406 1418 4444 1458
rect 4484 1418 4520 1458
rect 4406 1368 4520 1418
rect 5848 1558 5960 1608
rect 5848 1518 5884 1558
rect 5924 1518 5960 1558
rect 5848 1458 5960 1518
rect 5848 1418 5884 1458
rect 5924 1418 5960 1458
rect 5848 1368 5960 1418
rect 5990 1558 6104 1608
rect 5990 1518 6028 1558
rect 6068 1518 6104 1558
rect 5990 1458 6104 1518
rect 5990 1418 6028 1458
rect 6068 1418 6104 1458
rect 5990 1368 6104 1418
rect 6134 1558 6248 1608
rect 6134 1518 6172 1558
rect 6212 1518 6248 1558
rect 6134 1458 6248 1518
rect 6134 1418 6172 1458
rect 6212 1418 6248 1458
rect 6134 1368 6248 1418
rect 6424 1558 6536 1608
rect 6424 1518 6460 1558
rect 6500 1518 6536 1558
rect 6424 1458 6536 1518
rect 6424 1418 6460 1458
rect 6500 1418 6536 1458
rect 6424 1368 6536 1418
rect 6566 1558 6680 1608
rect 6566 1518 6604 1558
rect 6644 1518 6680 1558
rect 6566 1458 6680 1518
rect 6566 1418 6604 1458
rect 6644 1418 6680 1458
rect 6566 1368 6680 1418
rect 6710 1558 6824 1608
rect 6710 1518 6748 1558
rect 6788 1518 6824 1558
rect 6710 1458 6824 1518
rect 6710 1418 6748 1458
rect 6788 1418 6824 1458
rect 6710 1368 6824 1418
rect 7000 1558 7112 1608
rect 7000 1518 7036 1558
rect 7076 1518 7112 1558
rect 7000 1458 7112 1518
rect 7000 1418 7036 1458
rect 7076 1418 7112 1458
rect 7000 1368 7112 1418
rect 7142 1558 7256 1608
rect 7142 1518 7180 1558
rect 7220 1518 7256 1558
rect 7142 1458 7256 1518
rect 7142 1418 7180 1458
rect 7220 1418 7256 1458
rect 7142 1368 7256 1418
rect 7286 1558 7400 1608
rect 7286 1518 7324 1558
rect 7364 1518 7400 1558
rect 7286 1458 7400 1518
rect 7286 1418 7324 1458
rect 7364 1418 7400 1458
rect 7286 1368 7400 1418
rect 7576 1558 7688 1608
rect 7576 1518 7612 1558
rect 7652 1518 7688 1558
rect 7576 1458 7688 1518
rect 7576 1418 7612 1458
rect 7652 1418 7688 1458
rect 7576 1368 7688 1418
rect 7718 1558 7832 1608
rect 7718 1518 7756 1558
rect 7796 1518 7832 1558
rect 7718 1458 7832 1518
rect 7718 1418 7756 1458
rect 7796 1418 7832 1458
rect 7718 1368 7832 1418
rect 7862 1558 7976 1608
rect 7862 1518 7900 1558
rect 7940 1518 7976 1558
rect 7862 1458 7976 1518
rect 7862 1418 7900 1458
rect 7940 1418 7976 1458
rect 7862 1368 7976 1418
rect 8152 1558 8264 1608
rect 8152 1518 8188 1558
rect 8228 1518 8264 1558
rect 8152 1458 8264 1518
rect 8152 1418 8188 1458
rect 8228 1418 8264 1458
rect 8152 1368 8264 1418
rect 8294 1558 8408 1608
rect 8294 1518 8332 1558
rect 8372 1518 8408 1558
rect 8294 1458 8408 1518
rect 8294 1418 8332 1458
rect 8372 1418 8408 1458
rect 8294 1368 8408 1418
rect 8438 1558 8552 1608
rect 8438 1518 8476 1558
rect 8516 1518 8552 1558
rect 8438 1458 8552 1518
rect 8438 1418 8476 1458
rect 8516 1418 8552 1458
rect 8438 1368 8552 1418
rect 9304 1558 9416 1608
rect 9304 1518 9340 1558
rect 9380 1518 9416 1558
rect 9304 1458 9416 1518
rect 9304 1418 9340 1458
rect 9380 1418 9416 1458
rect 9304 1368 9416 1418
rect 9446 1558 9560 1608
rect 9446 1518 9484 1558
rect 9524 1518 9560 1558
rect 9446 1458 9560 1518
rect 9446 1418 9484 1458
rect 9524 1418 9560 1458
rect 9446 1368 9560 1418
rect 9590 1558 9704 1608
rect 9590 1518 9628 1558
rect 9668 1518 9704 1558
rect 9590 1458 9704 1518
rect 9590 1418 9628 1458
rect 9668 1418 9704 1458
rect 9590 1368 9704 1418
rect 9880 1558 9992 1608
rect 9880 1518 9916 1558
rect 9956 1518 9992 1558
rect 9880 1458 9992 1518
rect 9880 1418 9916 1458
rect 9956 1418 9992 1458
rect 9880 1368 9992 1418
rect 10022 1558 10136 1608
rect 10022 1518 10060 1558
rect 10100 1518 10136 1558
rect 10022 1458 10136 1518
rect 10022 1418 10060 1458
rect 10100 1418 10136 1458
rect 10022 1368 10136 1418
rect 10166 1558 10280 1608
rect 10166 1518 10204 1558
rect 10244 1518 10280 1558
rect 10166 1458 10280 1518
rect 10166 1418 10204 1458
rect 10244 1418 10280 1458
rect 10166 1368 10280 1418
rect 10456 1558 10568 1608
rect 10456 1518 10492 1558
rect 10532 1518 10568 1558
rect 10456 1458 10568 1518
rect 10456 1418 10492 1458
rect 10532 1418 10568 1458
rect 10456 1368 10568 1418
rect 10598 1558 10712 1608
rect 10598 1518 10636 1558
rect 10676 1518 10712 1558
rect 10598 1458 10712 1518
rect 10598 1418 10636 1458
rect 10676 1418 10712 1458
rect 10598 1368 10712 1418
rect 10742 1558 10856 1608
rect 10742 1518 10780 1558
rect 10820 1518 10856 1558
rect 10742 1458 10856 1518
rect 10742 1418 10780 1458
rect 10820 1418 10856 1458
rect 10742 1368 10856 1418
rect 11032 1558 11144 1608
rect 11032 1518 11068 1558
rect 11108 1518 11144 1558
rect 11032 1458 11144 1518
rect 11032 1418 11068 1458
rect 11108 1418 11144 1458
rect 11032 1368 11144 1418
rect 11174 1558 11288 1608
rect 11174 1518 11212 1558
rect 11252 1518 11288 1558
rect 11174 1458 11288 1518
rect 11174 1418 11212 1458
rect 11252 1418 11288 1458
rect 11174 1368 11288 1418
rect 11318 1558 11432 1608
rect 11318 1518 11356 1558
rect 11396 1518 11432 1558
rect 11318 1458 11432 1518
rect 11318 1418 11356 1458
rect 11396 1418 11432 1458
rect 11318 1368 11432 1418
rect 11896 1558 12008 1608
rect 11896 1518 11932 1558
rect 11972 1518 12008 1558
rect 11896 1458 12008 1518
rect 11896 1418 11932 1458
rect 11972 1418 12008 1458
rect 11896 1368 12008 1418
rect 12038 1558 12152 1608
rect 12038 1518 12076 1558
rect 12116 1518 12152 1558
rect 12038 1458 12152 1518
rect 12038 1418 12076 1458
rect 12116 1418 12152 1458
rect 12038 1368 12152 1418
rect 12182 1558 12296 1608
rect 12182 1518 12220 1558
rect 12260 1518 12296 1558
rect 12182 1458 12296 1518
rect 12182 1418 12220 1458
rect 12260 1418 12296 1458
rect 12182 1368 12296 1418
rect 12472 1558 12584 1608
rect 12472 1518 12508 1558
rect 12548 1518 12584 1558
rect 12472 1458 12584 1518
rect 12472 1418 12508 1458
rect 12548 1418 12584 1458
rect 12472 1368 12584 1418
rect 12614 1558 12728 1608
rect 12614 1518 12652 1558
rect 12692 1518 12728 1558
rect 12614 1458 12728 1518
rect 12614 1418 12652 1458
rect 12692 1418 12728 1458
rect 12614 1368 12728 1418
rect 12758 1558 12872 1608
rect 12758 1518 12796 1558
rect 12836 1518 12872 1558
rect 12758 1458 12872 1518
rect 12758 1418 12796 1458
rect 12836 1418 12872 1458
rect 12758 1368 12872 1418
rect 13048 1558 13160 1608
rect 13048 1518 13084 1558
rect 13124 1518 13160 1558
rect 13048 1458 13160 1518
rect 13048 1418 13084 1458
rect 13124 1418 13160 1458
rect 13048 1368 13160 1418
rect 13190 1558 13304 1608
rect 13190 1518 13228 1558
rect 13268 1518 13304 1558
rect 13190 1458 13304 1518
rect 13190 1418 13228 1458
rect 13268 1418 13304 1458
rect 13190 1368 13304 1418
rect 13334 1558 13448 1608
rect 13334 1518 13372 1558
rect 13412 1518 13448 1558
rect 13334 1458 13448 1518
rect 13334 1418 13372 1458
rect 13412 1418 13448 1458
rect 13334 1368 13448 1418
rect 13624 1558 13736 1608
rect 13624 1518 13660 1558
rect 13700 1518 13736 1558
rect 13624 1458 13736 1518
rect 13624 1418 13660 1458
rect 13700 1418 13736 1458
rect 13624 1368 13736 1418
rect 13766 1558 13880 1608
rect 13766 1518 13804 1558
rect 13844 1518 13880 1558
rect 13766 1458 13880 1518
rect 13766 1418 13804 1458
rect 13844 1418 13880 1458
rect 13766 1368 13880 1418
rect 13910 1558 14024 1608
rect 13910 1518 13948 1558
rect 13988 1518 14024 1558
rect 13910 1458 14024 1518
rect 13910 1418 13948 1458
rect 13988 1418 14024 1458
rect 13910 1368 14024 1418
rect 14776 1558 14888 1608
rect 14776 1518 14812 1558
rect 14852 1518 14888 1558
rect 14776 1458 14888 1518
rect 14776 1418 14812 1458
rect 14852 1418 14888 1458
rect 14776 1368 14888 1418
rect 14918 1558 15032 1608
rect 14918 1518 14956 1558
rect 14996 1518 15032 1558
rect 14918 1458 15032 1518
rect 14918 1418 14956 1458
rect 14996 1418 15032 1458
rect 14918 1368 15032 1418
rect 15062 1558 15176 1608
rect 15062 1518 15100 1558
rect 15140 1518 15176 1558
rect 15062 1458 15176 1518
rect 15062 1418 15100 1458
rect 15140 1418 15176 1458
rect 15062 1368 15176 1418
rect 15352 1558 15466 1608
rect 15352 1518 15388 1558
rect 15428 1518 15466 1558
rect 15352 1458 15466 1518
rect 15352 1418 15388 1458
rect 15428 1418 15466 1458
rect 15352 1368 15466 1418
rect 15496 1558 15610 1608
rect 15496 1518 15532 1558
rect 15572 1518 15610 1558
rect 15496 1458 15610 1518
rect 15496 1418 15532 1458
rect 15572 1418 15610 1458
rect 15496 1368 15610 1418
rect 15640 1558 15752 1608
rect 15640 1518 15676 1558
rect 15716 1518 15752 1558
rect 15640 1458 15752 1518
rect 15640 1418 15676 1458
rect 15716 1418 15752 1458
rect 15640 1368 15752 1418
rect 15928 1558 16040 1608
rect 15928 1518 15964 1558
rect 16004 1518 16040 1558
rect 15928 1458 16040 1518
rect 15928 1418 15964 1458
rect 16004 1418 16040 1458
rect 15928 1368 16040 1418
rect 16070 1558 16184 1608
rect 16070 1518 16108 1558
rect 16148 1518 16184 1558
rect 16070 1458 16184 1518
rect 16070 1418 16108 1458
rect 16148 1418 16184 1458
rect 16070 1368 16184 1418
rect 16214 1558 16328 1608
rect 16214 1518 16252 1558
rect 16292 1518 16328 1558
rect 16214 1458 16328 1518
rect 16214 1418 16252 1458
rect 16292 1418 16328 1458
rect 16214 1368 16328 1418
rect 16358 1558 16472 1608
rect 16358 1518 16396 1558
rect 16436 1518 16472 1558
rect 16358 1458 16472 1518
rect 16358 1418 16396 1458
rect 16436 1418 16472 1458
rect 16358 1368 16472 1418
rect 16502 1558 16616 1608
rect 16502 1518 16540 1558
rect 16580 1518 16616 1558
rect 16502 1458 16616 1518
rect 16502 1418 16540 1458
rect 16580 1418 16616 1458
rect 16502 1368 16616 1418
rect 17368 1558 17480 1608
rect 17368 1518 17404 1558
rect 17444 1518 17480 1558
rect 17368 1458 17480 1518
rect 17368 1418 17404 1458
rect 17444 1418 17480 1458
rect 17368 1368 17480 1418
rect 17510 1558 17624 1608
rect 17510 1518 17548 1558
rect 17588 1518 17624 1558
rect 17510 1458 17624 1518
rect 17510 1418 17548 1458
rect 17588 1418 17624 1458
rect 17510 1368 17624 1418
rect 17654 1558 17768 1608
rect 17654 1518 17692 1558
rect 17732 1518 17768 1558
rect 17654 1458 17768 1518
rect 17654 1418 17692 1458
rect 17732 1418 17768 1458
rect 17654 1368 17768 1418
rect 17798 1558 17912 1608
rect 17798 1518 17836 1558
rect 17876 1518 17912 1558
rect 17798 1458 17912 1518
rect 17798 1418 17836 1458
rect 17876 1418 17912 1458
rect 17798 1368 17912 1418
rect 17942 1558 18056 1608
rect 17942 1518 17980 1558
rect 18020 1518 18056 1558
rect 17942 1458 18056 1518
rect 17942 1418 17980 1458
rect 18020 1418 18056 1458
rect 17942 1368 18056 1418
rect 18086 1558 18200 1608
rect 18086 1518 18124 1558
rect 18164 1518 18200 1558
rect 18086 1458 18200 1518
rect 18086 1418 18124 1458
rect 18164 1418 18200 1458
rect 18086 1368 18200 1418
rect 18230 1558 18344 1608
rect 18230 1518 18268 1558
rect 18308 1518 18344 1558
rect 18230 1458 18344 1518
rect 18230 1418 18268 1458
rect 18308 1418 18344 1458
rect 18230 1368 18344 1418
rect 18374 1558 18488 1608
rect 18374 1518 18412 1558
rect 18452 1518 18488 1558
rect 18374 1458 18488 1518
rect 18374 1418 18412 1458
rect 18452 1418 18488 1458
rect 18374 1368 18488 1418
rect 18518 1558 18632 1608
rect 18518 1518 18556 1558
rect 18596 1518 18632 1558
rect 18518 1458 18632 1518
rect 18518 1418 18556 1458
rect 18596 1418 18632 1458
rect 18518 1368 18632 1418
rect 18662 1558 18776 1608
rect 18662 1518 18700 1558
rect 18740 1518 18776 1558
rect 18662 1458 18776 1518
rect 18662 1418 18700 1458
rect 18740 1418 18776 1458
rect 18662 1368 18776 1418
rect 18806 1558 18920 1608
rect 18806 1518 18844 1558
rect 18884 1518 18920 1558
rect 18806 1458 18920 1518
rect 18806 1418 18844 1458
rect 18884 1418 18920 1458
rect 18806 1368 18920 1418
rect 18950 1558 19064 1608
rect 18950 1518 18988 1558
rect 19028 1518 19064 1558
rect 18950 1458 19064 1518
rect 18950 1418 18988 1458
rect 19028 1418 19064 1458
rect 18950 1368 19064 1418
rect 19094 1558 19208 1608
rect 19094 1518 19132 1558
rect 19172 1518 19208 1558
rect 19094 1458 19208 1518
rect 19094 1418 19132 1458
rect 19172 1418 19208 1458
rect 19094 1368 19208 1418
rect 19238 1558 19352 1608
rect 19238 1518 19276 1558
rect 19316 1518 19352 1558
rect 19238 1458 19352 1518
rect 19238 1418 19276 1458
rect 19316 1418 19352 1458
rect 19238 1368 19352 1418
rect 19382 1558 19496 1608
rect 19382 1518 19420 1558
rect 19460 1518 19496 1558
rect 19382 1458 19496 1518
rect 19382 1418 19420 1458
rect 19460 1418 19496 1458
rect 19382 1368 19496 1418
rect 19526 1558 19640 1608
rect 19526 1518 19564 1558
rect 19604 1518 19640 1558
rect 19526 1458 19640 1518
rect 19526 1418 19564 1458
rect 19604 1418 19640 1458
rect 19526 1368 19640 1418
rect 19670 1558 19784 1608
rect 19670 1518 19708 1558
rect 19748 1518 19784 1558
rect 19670 1458 19784 1518
rect 19670 1418 19708 1458
rect 19748 1418 19784 1458
rect 19670 1368 19784 1418
rect 19814 1558 19928 1608
rect 19814 1518 19852 1558
rect 19892 1518 19928 1558
rect 19814 1458 19928 1518
rect 19814 1418 19852 1458
rect 19892 1418 19928 1458
rect 19814 1368 19928 1418
rect 19958 1558 20072 1608
rect 19958 1518 19996 1558
rect 20036 1518 20072 1558
rect 19958 1458 20072 1518
rect 19958 1418 19996 1458
rect 20036 1418 20072 1458
rect 19958 1368 20072 1418
rect 20102 1558 20216 1608
rect 20102 1518 20140 1558
rect 20180 1518 20216 1558
rect 20102 1458 20216 1518
rect 20102 1418 20140 1458
rect 20180 1418 20216 1458
rect 20102 1368 20216 1418
rect 20246 1558 20360 1608
rect 20246 1518 20284 1558
rect 20324 1518 20360 1558
rect 20246 1458 20360 1518
rect 20246 1418 20284 1458
rect 20324 1418 20360 1458
rect 20246 1368 20360 1418
rect 20390 1558 20504 1608
rect 20390 1518 20428 1558
rect 20468 1518 20504 1558
rect 20390 1458 20504 1518
rect 20390 1418 20428 1458
rect 20468 1418 20504 1458
rect 20390 1368 20504 1418
rect 20534 1558 20648 1608
rect 20534 1518 20572 1558
rect 20612 1518 20648 1558
rect 20534 1458 20648 1518
rect 20534 1418 20572 1458
rect 20612 1418 20648 1458
rect 20534 1368 20648 1418
rect 20678 1558 20792 1608
rect 20678 1518 20716 1558
rect 20756 1518 20792 1558
rect 20678 1458 20792 1518
rect 20678 1418 20716 1458
rect 20756 1418 20792 1458
rect 20678 1368 20792 1418
rect 20822 1558 20936 1608
rect 20822 1518 20860 1558
rect 20900 1518 20936 1558
rect 20822 1458 20936 1518
rect 20822 1418 20860 1458
rect 20900 1418 20936 1458
rect 20822 1368 20936 1418
<< pdiff >>
rect 664 3794 778 3864
rect 664 3754 700 3794
rect 740 3754 778 3794
rect 664 3694 778 3754
rect 664 3654 700 3694
rect 740 3654 778 3694
rect 664 3594 778 3654
rect 664 3554 700 3594
rect 740 3554 778 3594
rect 664 3494 778 3554
rect 664 3454 700 3494
rect 740 3454 778 3494
rect 664 3384 778 3454
rect 808 3794 922 3864
rect 808 3754 844 3794
rect 884 3754 922 3794
rect 808 3694 922 3754
rect 808 3654 844 3694
rect 884 3654 922 3694
rect 808 3594 922 3654
rect 808 3554 844 3594
rect 884 3554 922 3594
rect 808 3494 922 3554
rect 808 3454 844 3494
rect 884 3454 922 3494
rect 808 3384 922 3454
rect 952 3794 1064 3864
rect 952 3754 988 3794
rect 1028 3754 1064 3794
rect 952 3694 1064 3754
rect 952 3654 988 3694
rect 1028 3654 1064 3694
rect 952 3594 1064 3654
rect 952 3554 988 3594
rect 1028 3554 1064 3594
rect 952 3494 1064 3554
rect 952 3454 988 3494
rect 1028 3454 1064 3494
rect 952 3384 1064 3454
rect 1240 3794 1354 3864
rect 1240 3754 1276 3794
rect 1316 3754 1354 3794
rect 1240 3694 1354 3754
rect 1240 3654 1276 3694
rect 1316 3654 1354 3694
rect 1240 3594 1354 3654
rect 1240 3554 1276 3594
rect 1316 3554 1354 3594
rect 1240 3494 1354 3554
rect 1240 3454 1276 3494
rect 1316 3454 1354 3494
rect 1240 3384 1354 3454
rect 1384 3794 1498 3864
rect 1384 3754 1420 3794
rect 1460 3754 1498 3794
rect 1384 3694 1498 3754
rect 1384 3654 1420 3694
rect 1460 3654 1498 3694
rect 1384 3594 1498 3654
rect 1384 3554 1420 3594
rect 1460 3554 1498 3594
rect 1384 3494 1498 3554
rect 1384 3454 1420 3494
rect 1460 3454 1498 3494
rect 1384 3384 1498 3454
rect 1528 3794 1640 3864
rect 1528 3754 1564 3794
rect 1604 3754 1640 3794
rect 1528 3694 1640 3754
rect 1528 3654 1564 3694
rect 1604 3654 1640 3694
rect 1528 3594 1640 3654
rect 1528 3554 1564 3594
rect 1604 3554 1640 3594
rect 1528 3494 1640 3554
rect 1528 3454 1564 3494
rect 1604 3454 1640 3494
rect 1528 3384 1640 3454
rect 1816 3794 1930 3864
rect 1816 3754 1852 3794
rect 1892 3754 1930 3794
rect 1816 3694 1930 3754
rect 1816 3654 1852 3694
rect 1892 3654 1930 3694
rect 1816 3594 1930 3654
rect 1816 3554 1852 3594
rect 1892 3554 1930 3594
rect 1816 3494 1930 3554
rect 1816 3454 1852 3494
rect 1892 3454 1930 3494
rect 1816 3384 1930 3454
rect 1960 3794 2074 3864
rect 1960 3754 1996 3794
rect 2036 3754 2074 3794
rect 1960 3694 2074 3754
rect 1960 3654 1996 3694
rect 2036 3654 2074 3694
rect 1960 3594 2074 3654
rect 1960 3554 1996 3594
rect 2036 3554 2074 3594
rect 1960 3494 2074 3554
rect 1960 3454 1996 3494
rect 2036 3454 2074 3494
rect 1960 3384 2074 3454
rect 2104 3794 2216 3864
rect 2104 3754 2140 3794
rect 2180 3754 2216 3794
rect 2104 3694 2216 3754
rect 2104 3654 2140 3694
rect 2180 3654 2216 3694
rect 2104 3594 2216 3654
rect 2104 3554 2140 3594
rect 2180 3554 2216 3594
rect 2104 3494 2216 3554
rect 2104 3454 2140 3494
rect 2180 3454 2216 3494
rect 2104 3384 2216 3454
rect 2392 3794 2506 3864
rect 2392 3754 2428 3794
rect 2468 3754 2506 3794
rect 2392 3694 2506 3754
rect 2392 3654 2428 3694
rect 2468 3654 2506 3694
rect 2392 3594 2506 3654
rect 2392 3554 2428 3594
rect 2468 3554 2506 3594
rect 2392 3494 2506 3554
rect 2392 3454 2428 3494
rect 2468 3454 2506 3494
rect 2392 3384 2506 3454
rect 2536 3794 2650 3864
rect 2536 3754 2572 3794
rect 2612 3754 2650 3794
rect 2536 3694 2650 3754
rect 2536 3654 2572 3694
rect 2612 3654 2650 3694
rect 2536 3594 2650 3654
rect 2536 3554 2572 3594
rect 2612 3554 2650 3594
rect 2536 3494 2650 3554
rect 2536 3454 2572 3494
rect 2612 3454 2650 3494
rect 2536 3384 2650 3454
rect 2680 3794 2792 3864
rect 2680 3754 2716 3794
rect 2756 3754 2792 3794
rect 2680 3694 2792 3754
rect 2680 3654 2716 3694
rect 2756 3654 2792 3694
rect 2680 3594 2792 3654
rect 2680 3554 2716 3594
rect 2756 3554 2792 3594
rect 2680 3494 2792 3554
rect 2680 3454 2716 3494
rect 2756 3454 2792 3494
rect 2680 3384 2792 3454
rect 2968 3794 3080 3864
rect 2968 3754 3004 3794
rect 3044 3754 3080 3794
rect 2968 3694 3080 3754
rect 2968 3654 3004 3694
rect 3044 3654 3080 3694
rect 2968 3594 3080 3654
rect 2968 3554 3004 3594
rect 3044 3554 3080 3594
rect 2968 3494 3080 3554
rect 2968 3454 3004 3494
rect 3044 3454 3080 3494
rect 2968 3384 3080 3454
rect 3110 3794 3224 3864
rect 3110 3754 3148 3794
rect 3188 3754 3224 3794
rect 3110 3694 3224 3754
rect 3110 3654 3148 3694
rect 3188 3654 3224 3694
rect 3110 3594 3224 3654
rect 3110 3554 3148 3594
rect 3188 3554 3224 3594
rect 3110 3494 3224 3554
rect 3110 3454 3148 3494
rect 3188 3454 3224 3494
rect 3110 3384 3224 3454
rect 3254 3794 3368 3864
rect 3254 3754 3292 3794
rect 3332 3754 3368 3794
rect 3254 3694 3368 3754
rect 4120 3794 4232 3864
rect 4120 3754 4156 3794
rect 4196 3754 4232 3794
rect 3254 3654 3292 3694
rect 3332 3654 3368 3694
rect 3254 3594 3368 3654
rect 3254 3554 3292 3594
rect 3332 3554 3368 3594
rect 3254 3494 3368 3554
rect 4120 3694 4232 3754
rect 4120 3654 4156 3694
rect 4196 3654 4232 3694
rect 4120 3594 4232 3654
rect 4120 3554 4156 3594
rect 4196 3554 4232 3594
rect 3254 3454 3292 3494
rect 3332 3454 3368 3494
rect 3254 3384 3368 3454
rect 4120 3494 4232 3554
rect 4120 3454 4156 3494
rect 4196 3454 4232 3494
rect 4120 3384 4232 3454
rect 4262 3794 4376 3864
rect 4262 3754 4300 3794
rect 4340 3754 4376 3794
rect 4262 3694 4376 3754
rect 4262 3654 4300 3694
rect 4340 3654 4376 3694
rect 4262 3594 4376 3654
rect 4262 3554 4300 3594
rect 4340 3554 4376 3594
rect 4262 3494 4376 3554
rect 4262 3454 4300 3494
rect 4340 3454 4376 3494
rect 4262 3384 4376 3454
rect 4406 3794 4520 3864
rect 4406 3754 4444 3794
rect 4484 3754 4520 3794
rect 4406 3694 4520 3754
rect 4406 3654 4444 3694
rect 4484 3654 4520 3694
rect 4406 3594 4520 3654
rect 4406 3554 4444 3594
rect 4484 3554 4520 3594
rect 4406 3494 4520 3554
rect 4406 3454 4444 3494
rect 4484 3454 4520 3494
rect 4406 3384 4520 3454
rect 4696 3794 4808 3864
rect 4696 3754 4732 3794
rect 4772 3754 4808 3794
rect 4696 3694 4808 3754
rect 4696 3654 4732 3694
rect 4772 3654 4808 3694
rect 4696 3594 4808 3654
rect 4696 3554 4732 3594
rect 4772 3554 4808 3594
rect 4696 3494 4808 3554
rect 4696 3454 4732 3494
rect 4772 3454 4808 3494
rect 4696 3384 4808 3454
rect 4838 3794 4952 3864
rect 4838 3754 4876 3794
rect 4916 3754 4952 3794
rect 4838 3694 4952 3754
rect 4838 3654 4876 3694
rect 4916 3654 4952 3694
rect 4838 3594 4952 3654
rect 4838 3554 4876 3594
rect 4916 3554 4952 3594
rect 4838 3494 4952 3554
rect 4838 3454 4876 3494
rect 4916 3454 4952 3494
rect 4838 3384 4952 3454
rect 4982 3794 5096 3864
rect 4982 3754 5020 3794
rect 5060 3754 5096 3794
rect 4982 3694 5096 3754
rect 4982 3654 5020 3694
rect 5060 3654 5096 3694
rect 4982 3594 5096 3654
rect 4982 3554 5020 3594
rect 5060 3554 5096 3594
rect 4982 3494 5096 3554
rect 4982 3454 5020 3494
rect 5060 3454 5096 3494
rect 4982 3384 5096 3454
rect 5272 3794 5384 3864
rect 5272 3754 5308 3794
rect 5348 3754 5384 3794
rect 5272 3694 5384 3754
rect 5272 3654 5308 3694
rect 5348 3654 5384 3694
rect 5272 3594 5384 3654
rect 5272 3554 5308 3594
rect 5348 3554 5384 3594
rect 5272 3494 5384 3554
rect 5272 3454 5308 3494
rect 5348 3454 5384 3494
rect 5272 3384 5384 3454
rect 5414 3794 5528 3864
rect 5414 3754 5452 3794
rect 5492 3754 5528 3794
rect 5414 3694 5528 3754
rect 5414 3654 5452 3694
rect 5492 3654 5528 3694
rect 5414 3594 5528 3654
rect 5414 3554 5452 3594
rect 5492 3554 5528 3594
rect 5414 3494 5528 3554
rect 5414 3454 5452 3494
rect 5492 3454 5528 3494
rect 5414 3384 5528 3454
rect 5558 3794 5672 3864
rect 5558 3754 5596 3794
rect 5636 3754 5672 3794
rect 5558 3694 5672 3754
rect 5558 3654 5596 3694
rect 5636 3654 5672 3694
rect 5558 3594 5672 3654
rect 5558 3554 5596 3594
rect 5636 3554 5672 3594
rect 5558 3494 5672 3554
rect 5558 3454 5596 3494
rect 5636 3454 5672 3494
rect 5558 3384 5672 3454
rect 5848 3794 5960 3864
rect 5848 3754 5884 3794
rect 5924 3754 5960 3794
rect 5848 3694 5960 3754
rect 5848 3654 5884 3694
rect 5924 3654 5960 3694
rect 5848 3594 5960 3654
rect 5848 3554 5884 3594
rect 5924 3554 5960 3594
rect 5848 3494 5960 3554
rect 5848 3454 5884 3494
rect 5924 3454 5960 3494
rect 5848 3384 5960 3454
rect 5990 3794 6104 3864
rect 5990 3754 6028 3794
rect 6068 3754 6104 3794
rect 5990 3694 6104 3754
rect 5990 3654 6028 3694
rect 6068 3654 6104 3694
rect 5990 3594 6104 3654
rect 5990 3554 6028 3594
rect 6068 3554 6104 3594
rect 5990 3494 6104 3554
rect 5990 3454 6028 3494
rect 6068 3454 6104 3494
rect 5990 3384 6104 3454
rect 6134 3794 6248 3864
rect 6134 3754 6172 3794
rect 6212 3754 6248 3794
rect 6134 3694 6248 3754
rect 6134 3654 6172 3694
rect 6212 3654 6248 3694
rect 6134 3594 6248 3654
rect 6134 3554 6172 3594
rect 6212 3554 6248 3594
rect 6134 3494 6248 3554
rect 6134 3454 6172 3494
rect 6212 3454 6248 3494
rect 6134 3384 6248 3454
rect 6424 3794 6536 3864
rect 6424 3754 6460 3794
rect 6500 3754 6536 3794
rect 6424 3694 6536 3754
rect 6424 3654 6460 3694
rect 6500 3654 6536 3694
rect 6424 3594 6536 3654
rect 6424 3554 6460 3594
rect 6500 3554 6536 3594
rect 6424 3494 6536 3554
rect 6424 3454 6460 3494
rect 6500 3454 6536 3494
rect 6424 3384 6536 3454
rect 6566 3794 6680 3864
rect 6566 3754 6604 3794
rect 6644 3754 6680 3794
rect 6566 3694 6680 3754
rect 6566 3654 6604 3694
rect 6644 3654 6680 3694
rect 6566 3594 6680 3654
rect 6566 3554 6604 3594
rect 6644 3554 6680 3594
rect 6566 3494 6680 3554
rect 6566 3454 6604 3494
rect 6644 3454 6680 3494
rect 6566 3384 6680 3454
rect 6710 3794 6824 3864
rect 6710 3754 6748 3794
rect 6788 3754 6824 3794
rect 6710 3694 6824 3754
rect 7576 3794 7688 3864
rect 7576 3754 7612 3794
rect 7652 3754 7688 3794
rect 6710 3654 6748 3694
rect 6788 3654 6824 3694
rect 6710 3594 6824 3654
rect 6710 3554 6748 3594
rect 6788 3554 6824 3594
rect 6710 3494 6824 3554
rect 7576 3694 7688 3754
rect 7576 3654 7612 3694
rect 7652 3654 7688 3694
rect 7576 3594 7688 3654
rect 7576 3554 7612 3594
rect 7652 3554 7688 3594
rect 6710 3454 6748 3494
rect 6788 3454 6824 3494
rect 6710 3384 6824 3454
rect 7576 3494 7688 3554
rect 7576 3454 7612 3494
rect 7652 3454 7688 3494
rect 7576 3384 7688 3454
rect 7718 3794 7832 3864
rect 7718 3754 7756 3794
rect 7796 3754 7832 3794
rect 7718 3694 7832 3754
rect 7718 3654 7756 3694
rect 7796 3654 7832 3694
rect 7718 3594 7832 3654
rect 7718 3554 7756 3594
rect 7796 3554 7832 3594
rect 7718 3494 7832 3554
rect 7718 3454 7756 3494
rect 7796 3454 7832 3494
rect 7718 3384 7832 3454
rect 7862 3794 7976 3864
rect 7862 3754 7900 3794
rect 7940 3754 7976 3794
rect 7862 3694 7976 3754
rect 7862 3654 7900 3694
rect 7940 3654 7976 3694
rect 7862 3594 7976 3654
rect 7862 3554 7900 3594
rect 7940 3554 7976 3594
rect 7862 3494 7976 3554
rect 7862 3454 7900 3494
rect 7940 3454 7976 3494
rect 7862 3384 7976 3454
rect 8152 3794 8264 3864
rect 8152 3754 8188 3794
rect 8228 3754 8264 3794
rect 8152 3694 8264 3754
rect 8152 3654 8188 3694
rect 8228 3654 8264 3694
rect 8152 3594 8264 3654
rect 8152 3554 8188 3594
rect 8228 3554 8264 3594
rect 8152 3494 8264 3554
rect 8152 3454 8188 3494
rect 8228 3454 8264 3494
rect 8152 3384 8264 3454
rect 8294 3794 8408 3864
rect 8294 3754 8332 3794
rect 8372 3754 8408 3794
rect 8294 3694 8408 3754
rect 8294 3654 8332 3694
rect 8372 3654 8408 3694
rect 8294 3594 8408 3654
rect 8294 3554 8332 3594
rect 8372 3554 8408 3594
rect 8294 3494 8408 3554
rect 8294 3454 8332 3494
rect 8372 3454 8408 3494
rect 8294 3384 8408 3454
rect 8438 3794 8552 3864
rect 8438 3754 8476 3794
rect 8516 3754 8552 3794
rect 8438 3694 8552 3754
rect 8438 3654 8476 3694
rect 8516 3654 8552 3694
rect 8438 3594 8552 3654
rect 8438 3554 8476 3594
rect 8516 3554 8552 3594
rect 8438 3494 8552 3554
rect 8438 3454 8476 3494
rect 8516 3454 8552 3494
rect 8438 3384 8552 3454
rect 8728 3794 8840 3864
rect 8728 3754 8764 3794
rect 8804 3754 8840 3794
rect 8728 3694 8840 3754
rect 8728 3654 8764 3694
rect 8804 3654 8840 3694
rect 8728 3594 8840 3654
rect 8728 3554 8764 3594
rect 8804 3554 8840 3594
rect 8728 3494 8840 3554
rect 8728 3454 8764 3494
rect 8804 3454 8840 3494
rect 8728 3384 8840 3454
rect 8870 3794 8984 3864
rect 8870 3754 8908 3794
rect 8948 3754 8984 3794
rect 8870 3694 8984 3754
rect 8870 3654 8908 3694
rect 8948 3654 8984 3694
rect 8870 3594 8984 3654
rect 8870 3554 8908 3594
rect 8948 3554 8984 3594
rect 8870 3494 8984 3554
rect 8870 3454 8908 3494
rect 8948 3454 8984 3494
rect 8870 3384 8984 3454
rect 9014 3794 9128 3864
rect 9014 3754 9052 3794
rect 9092 3754 9128 3794
rect 9014 3694 9128 3754
rect 9014 3654 9052 3694
rect 9092 3654 9128 3694
rect 9014 3594 9128 3654
rect 9014 3554 9052 3594
rect 9092 3554 9128 3594
rect 9014 3494 9128 3554
rect 9014 3454 9052 3494
rect 9092 3454 9128 3494
rect 9014 3384 9128 3454
rect 9304 3794 9416 3864
rect 9304 3754 9340 3794
rect 9380 3754 9416 3794
rect 9304 3694 9416 3754
rect 9304 3654 9340 3694
rect 9380 3654 9416 3694
rect 9304 3594 9416 3654
rect 9304 3554 9340 3594
rect 9380 3554 9416 3594
rect 9304 3494 9416 3554
rect 9304 3454 9340 3494
rect 9380 3454 9416 3494
rect 9304 3384 9416 3454
rect 9446 3794 9560 3864
rect 9446 3754 9484 3794
rect 9524 3754 9560 3794
rect 9446 3694 9560 3754
rect 9446 3654 9484 3694
rect 9524 3654 9560 3694
rect 9446 3594 9560 3654
rect 9446 3554 9484 3594
rect 9524 3554 9560 3594
rect 9446 3494 9560 3554
rect 9446 3454 9484 3494
rect 9524 3454 9560 3494
rect 9446 3384 9560 3454
rect 9590 3794 9704 3864
rect 9590 3754 9628 3794
rect 9668 3754 9704 3794
rect 9590 3694 9704 3754
rect 9590 3654 9628 3694
rect 9668 3654 9704 3694
rect 9590 3594 9704 3654
rect 9590 3554 9628 3594
rect 9668 3554 9704 3594
rect 9590 3494 9704 3554
rect 9590 3454 9628 3494
rect 9668 3454 9704 3494
rect 9590 3384 9704 3454
rect 10168 3794 10280 3864
rect 10168 3754 10204 3794
rect 10244 3754 10280 3794
rect 10168 3694 10280 3754
rect 10168 3654 10204 3694
rect 10244 3654 10280 3694
rect 10168 3594 10280 3654
rect 10168 3554 10204 3594
rect 10244 3554 10280 3594
rect 10168 3494 10280 3554
rect 10168 3454 10204 3494
rect 10244 3454 10280 3494
rect 10168 3384 10280 3454
rect 10310 3794 10424 3864
rect 10310 3754 10348 3794
rect 10388 3754 10424 3794
rect 10310 3694 10424 3754
rect 10310 3654 10348 3694
rect 10388 3654 10424 3694
rect 10310 3594 10424 3654
rect 10310 3554 10348 3594
rect 10388 3554 10424 3594
rect 10310 3494 10424 3554
rect 10310 3454 10348 3494
rect 10388 3454 10424 3494
rect 10310 3384 10424 3454
rect 10454 3794 10568 3864
rect 10454 3754 10492 3794
rect 10532 3754 10568 3794
rect 10454 3694 10568 3754
rect 10454 3654 10492 3694
rect 10532 3654 10568 3694
rect 10454 3594 10568 3654
rect 10454 3554 10492 3594
rect 10532 3554 10568 3594
rect 10454 3494 10568 3554
rect 10454 3454 10492 3494
rect 10532 3454 10568 3494
rect 10454 3384 10568 3454
rect 10744 3794 10856 3864
rect 10744 3754 10780 3794
rect 10820 3754 10856 3794
rect 10744 3694 10856 3754
rect 10744 3654 10780 3694
rect 10820 3654 10856 3694
rect 10744 3594 10856 3654
rect 10744 3554 10780 3594
rect 10820 3554 10856 3594
rect 10744 3494 10856 3554
rect 10744 3454 10780 3494
rect 10820 3454 10856 3494
rect 10744 3384 10856 3454
rect 10886 3794 11000 3864
rect 10886 3754 10924 3794
rect 10964 3754 11000 3794
rect 10886 3694 11000 3754
rect 10886 3654 10924 3694
rect 10964 3654 11000 3694
rect 10886 3594 11000 3654
rect 10886 3554 10924 3594
rect 10964 3554 11000 3594
rect 10886 3494 11000 3554
rect 10886 3454 10924 3494
rect 10964 3454 11000 3494
rect 10886 3384 11000 3454
rect 11030 3794 11144 3864
rect 11030 3754 11068 3794
rect 11108 3754 11144 3794
rect 11030 3694 11144 3754
rect 11896 3794 12008 3864
rect 11896 3754 11932 3794
rect 11972 3754 12008 3794
rect 11030 3654 11068 3694
rect 11108 3654 11144 3694
rect 11030 3594 11144 3654
rect 11030 3554 11068 3594
rect 11108 3554 11144 3594
rect 11030 3494 11144 3554
rect 11896 3694 12008 3754
rect 11896 3654 11932 3694
rect 11972 3654 12008 3694
rect 11896 3594 12008 3654
rect 11896 3554 11932 3594
rect 11972 3554 12008 3594
rect 11030 3454 11068 3494
rect 11108 3454 11144 3494
rect 11030 3384 11144 3454
rect 11896 3494 12008 3554
rect 11896 3454 11932 3494
rect 11972 3454 12008 3494
rect 11896 3384 12008 3454
rect 12038 3794 12152 3864
rect 12038 3754 12076 3794
rect 12116 3754 12152 3794
rect 12038 3694 12152 3754
rect 12038 3654 12076 3694
rect 12116 3654 12152 3694
rect 12038 3594 12152 3654
rect 12038 3554 12076 3594
rect 12116 3554 12152 3594
rect 12038 3494 12152 3554
rect 12038 3454 12076 3494
rect 12116 3454 12152 3494
rect 12038 3384 12152 3454
rect 12182 3794 12296 3864
rect 12182 3754 12220 3794
rect 12260 3754 12296 3794
rect 12182 3694 12296 3754
rect 12182 3654 12220 3694
rect 12260 3654 12296 3694
rect 12182 3594 12296 3654
rect 12182 3554 12220 3594
rect 12260 3554 12296 3594
rect 12182 3494 12296 3554
rect 12182 3454 12220 3494
rect 12260 3454 12296 3494
rect 12182 3384 12296 3454
rect 12472 3794 12584 3864
rect 12472 3754 12508 3794
rect 12548 3754 12584 3794
rect 12472 3694 12584 3754
rect 12472 3654 12508 3694
rect 12548 3654 12584 3694
rect 12472 3594 12584 3654
rect 12472 3554 12508 3594
rect 12548 3554 12584 3594
rect 12472 3494 12584 3554
rect 12472 3454 12508 3494
rect 12548 3454 12584 3494
rect 12472 3384 12584 3454
rect 12614 3794 12728 3864
rect 12614 3754 12652 3794
rect 12692 3754 12728 3794
rect 12614 3694 12728 3754
rect 12614 3654 12652 3694
rect 12692 3654 12728 3694
rect 12614 3594 12728 3654
rect 12614 3554 12652 3594
rect 12692 3554 12728 3594
rect 12614 3494 12728 3554
rect 12614 3454 12652 3494
rect 12692 3454 12728 3494
rect 12614 3384 12728 3454
rect 12758 3794 12872 3864
rect 12758 3754 12796 3794
rect 12836 3754 12872 3794
rect 12758 3694 12872 3754
rect 12758 3654 12796 3694
rect 12836 3654 12872 3694
rect 12758 3594 12872 3654
rect 12758 3554 12796 3594
rect 12836 3554 12872 3594
rect 12758 3494 12872 3554
rect 12758 3454 12796 3494
rect 12836 3454 12872 3494
rect 12758 3384 12872 3454
rect 13624 3794 13736 3864
rect 13624 3754 13660 3794
rect 13700 3754 13736 3794
rect 13624 3694 13736 3754
rect 13624 3654 13660 3694
rect 13700 3654 13736 3694
rect 13624 3594 13736 3654
rect 13624 3554 13660 3594
rect 13700 3554 13736 3594
rect 13624 3494 13736 3554
rect 13624 3454 13660 3494
rect 13700 3454 13736 3494
rect 13624 3384 13736 3454
rect 13766 3794 13880 3864
rect 13766 3754 13804 3794
rect 13844 3754 13880 3794
rect 13766 3694 13880 3754
rect 13766 3654 13804 3694
rect 13844 3654 13880 3694
rect 13766 3594 13880 3654
rect 13766 3554 13804 3594
rect 13844 3554 13880 3594
rect 13766 3494 13880 3554
rect 13766 3454 13804 3494
rect 13844 3454 13880 3494
rect 13766 3384 13880 3454
rect 13910 3794 14024 3864
rect 13910 3754 13948 3794
rect 13988 3754 14024 3794
rect 13910 3694 14024 3754
rect 13910 3654 13948 3694
rect 13988 3654 14024 3694
rect 13910 3594 14024 3654
rect 13910 3554 13948 3594
rect 13988 3554 14024 3594
rect 13910 3494 14024 3554
rect 13910 3454 13948 3494
rect 13988 3454 14024 3494
rect 13910 3384 14024 3454
rect 14200 3794 14312 3864
rect 14200 3754 14236 3794
rect 14276 3754 14312 3794
rect 14200 3694 14312 3754
rect 14200 3654 14236 3694
rect 14276 3654 14312 3694
rect 14200 3594 14312 3654
rect 14200 3554 14236 3594
rect 14276 3554 14312 3594
rect 14200 3494 14312 3554
rect 14200 3454 14236 3494
rect 14276 3454 14312 3494
rect 14200 3384 14312 3454
rect 14342 3794 14456 3864
rect 14342 3754 14380 3794
rect 14420 3754 14456 3794
rect 14342 3694 14456 3754
rect 14342 3654 14380 3694
rect 14420 3654 14456 3694
rect 14342 3594 14456 3654
rect 14342 3554 14380 3594
rect 14420 3554 14456 3594
rect 14342 3494 14456 3554
rect 14342 3454 14380 3494
rect 14420 3454 14456 3494
rect 14342 3384 14456 3454
rect 14486 3794 14600 3864
rect 14486 3754 14524 3794
rect 14564 3754 14600 3794
rect 14486 3694 14600 3754
rect 14486 3654 14524 3694
rect 14564 3654 14600 3694
rect 14486 3594 14600 3654
rect 14486 3554 14524 3594
rect 14564 3554 14600 3594
rect 14486 3494 14600 3554
rect 14486 3454 14524 3494
rect 14564 3454 14600 3494
rect 14486 3384 14600 3454
rect 14776 3794 14888 3864
rect 14776 3754 14812 3794
rect 14852 3754 14888 3794
rect 14776 3694 14888 3754
rect 14776 3654 14812 3694
rect 14852 3654 14888 3694
rect 14776 3594 14888 3654
rect 14776 3554 14812 3594
rect 14852 3554 14888 3594
rect 14776 3494 14888 3554
rect 14776 3454 14812 3494
rect 14852 3454 14888 3494
rect 14776 3384 14888 3454
rect 14918 3794 15032 3864
rect 14918 3754 14956 3794
rect 14996 3754 15032 3794
rect 14918 3694 15032 3754
rect 14918 3654 14956 3694
rect 14996 3654 15032 3694
rect 14918 3594 15032 3654
rect 14918 3554 14956 3594
rect 14996 3554 15032 3594
rect 14918 3494 15032 3554
rect 14918 3454 14956 3494
rect 14996 3454 15032 3494
rect 14918 3384 15032 3454
rect 15062 3794 15176 3864
rect 15062 3754 15100 3794
rect 15140 3754 15176 3794
rect 15062 3694 15176 3754
rect 16504 3794 16618 3864
rect 16504 3754 16540 3794
rect 16580 3754 16618 3794
rect 15062 3654 15100 3694
rect 15140 3654 15176 3694
rect 15062 3594 15176 3654
rect 15062 3554 15100 3594
rect 15140 3554 15176 3594
rect 15062 3494 15176 3554
rect 16504 3694 16618 3754
rect 16504 3654 16540 3694
rect 16580 3654 16618 3694
rect 16504 3594 16618 3654
rect 16504 3554 16540 3594
rect 16580 3554 16618 3594
rect 15062 3454 15100 3494
rect 15140 3454 15176 3494
rect 15062 3384 15176 3454
rect 16504 3494 16618 3554
rect 16504 3454 16540 3494
rect 16580 3454 16618 3494
rect 16504 3384 16618 3454
rect 16648 3794 16762 3864
rect 16648 3754 16684 3794
rect 16724 3754 16762 3794
rect 16648 3694 16762 3754
rect 16648 3654 16684 3694
rect 16724 3654 16762 3694
rect 16648 3594 16762 3654
rect 16648 3554 16684 3594
rect 16724 3554 16762 3594
rect 16648 3494 16762 3554
rect 16648 3454 16684 3494
rect 16724 3454 16762 3494
rect 16648 3384 16762 3454
rect 16792 3794 16906 3864
rect 16792 3754 16828 3794
rect 16868 3754 16906 3794
rect 16792 3694 16906 3754
rect 16792 3654 16828 3694
rect 16868 3654 16906 3694
rect 16792 3594 16906 3654
rect 16792 3554 16828 3594
rect 16868 3554 16906 3594
rect 16792 3494 16906 3554
rect 16792 3454 16828 3494
rect 16868 3454 16906 3494
rect 16792 3384 16906 3454
rect 16936 3794 17050 3864
rect 16936 3754 16972 3794
rect 17012 3754 17050 3794
rect 16936 3694 17050 3754
rect 16936 3654 16972 3694
rect 17012 3654 17050 3694
rect 16936 3594 17050 3654
rect 16936 3554 16972 3594
rect 17012 3554 17050 3594
rect 16936 3494 17050 3554
rect 16936 3454 16972 3494
rect 17012 3454 17050 3494
rect 16936 3384 17050 3454
rect 17080 3794 17194 3864
rect 17080 3754 17116 3794
rect 17156 3754 17194 3794
rect 17080 3694 17194 3754
rect 17080 3654 17116 3694
rect 17156 3654 17194 3694
rect 17080 3594 17194 3654
rect 17080 3554 17116 3594
rect 17156 3554 17194 3594
rect 17080 3494 17194 3554
rect 17080 3454 17116 3494
rect 17156 3454 17194 3494
rect 17080 3384 17194 3454
rect 17224 3794 17338 3864
rect 17224 3754 17260 3794
rect 17300 3754 17338 3794
rect 17224 3694 17338 3754
rect 17224 3654 17260 3694
rect 17300 3654 17338 3694
rect 17224 3594 17338 3654
rect 17224 3554 17260 3594
rect 17300 3554 17338 3594
rect 17224 3494 17338 3554
rect 17224 3454 17260 3494
rect 17300 3454 17338 3494
rect 17224 3384 17338 3454
rect 17368 3794 17482 3864
rect 17368 3754 17404 3794
rect 17444 3754 17482 3794
rect 17368 3694 17482 3754
rect 17368 3654 17404 3694
rect 17444 3654 17482 3694
rect 17368 3594 17482 3654
rect 17368 3554 17404 3594
rect 17444 3554 17482 3594
rect 17368 3494 17482 3554
rect 17368 3454 17404 3494
rect 17444 3454 17482 3494
rect 17368 3384 17482 3454
rect 17512 3794 17626 3864
rect 17512 3754 17548 3794
rect 17588 3754 17626 3794
rect 17512 3694 17626 3754
rect 17512 3654 17548 3694
rect 17588 3654 17626 3694
rect 17512 3594 17626 3654
rect 17512 3554 17548 3594
rect 17588 3554 17626 3594
rect 17512 3494 17626 3554
rect 17512 3454 17548 3494
rect 17588 3454 17626 3494
rect 17512 3384 17626 3454
rect 17656 3794 17770 3864
rect 17656 3754 17692 3794
rect 17732 3754 17770 3794
rect 17656 3694 17770 3754
rect 17656 3654 17692 3694
rect 17732 3654 17770 3694
rect 17656 3594 17770 3654
rect 17656 3554 17692 3594
rect 17732 3554 17770 3594
rect 17656 3494 17770 3554
rect 17656 3454 17692 3494
rect 17732 3454 17770 3494
rect 17656 3384 17770 3454
rect 17800 3794 17914 3864
rect 17800 3754 17836 3794
rect 17876 3754 17914 3794
rect 17800 3694 17914 3754
rect 17800 3654 17836 3694
rect 17876 3654 17914 3694
rect 17800 3594 17914 3654
rect 17800 3554 17836 3594
rect 17876 3554 17914 3594
rect 17800 3494 17914 3554
rect 17800 3454 17836 3494
rect 17876 3454 17914 3494
rect 17800 3384 17914 3454
rect 17944 3794 18058 3864
rect 17944 3754 17980 3794
rect 18020 3754 18058 3794
rect 17944 3694 18058 3754
rect 17944 3654 17980 3694
rect 18020 3654 18058 3694
rect 17944 3594 18058 3654
rect 17944 3554 17980 3594
rect 18020 3554 18058 3594
rect 17944 3494 18058 3554
rect 17944 3454 17980 3494
rect 18020 3454 18058 3494
rect 17944 3384 18058 3454
rect 18088 3794 18202 3864
rect 18088 3754 18124 3794
rect 18164 3754 18202 3794
rect 18088 3694 18202 3754
rect 18088 3654 18124 3694
rect 18164 3654 18202 3694
rect 18088 3594 18202 3654
rect 18088 3554 18124 3594
rect 18164 3554 18202 3594
rect 18088 3494 18202 3554
rect 18088 3454 18124 3494
rect 18164 3454 18202 3494
rect 18088 3384 18202 3454
rect 18232 3794 18346 3864
rect 18232 3754 18268 3794
rect 18308 3754 18346 3794
rect 18232 3694 18346 3754
rect 18232 3654 18268 3694
rect 18308 3654 18346 3694
rect 18232 3594 18346 3654
rect 18232 3554 18268 3594
rect 18308 3554 18346 3594
rect 18232 3494 18346 3554
rect 18232 3454 18268 3494
rect 18308 3454 18346 3494
rect 18232 3384 18346 3454
rect 18376 3794 18490 3864
rect 18376 3754 18412 3794
rect 18452 3754 18490 3794
rect 18376 3694 18490 3754
rect 18376 3654 18412 3694
rect 18452 3654 18490 3694
rect 18376 3594 18490 3654
rect 18376 3554 18412 3594
rect 18452 3554 18490 3594
rect 18376 3494 18490 3554
rect 18376 3454 18412 3494
rect 18452 3454 18490 3494
rect 18376 3384 18490 3454
rect 18520 3794 18634 3864
rect 18520 3754 18556 3794
rect 18596 3754 18634 3794
rect 18520 3694 18634 3754
rect 18520 3654 18556 3694
rect 18596 3654 18634 3694
rect 18520 3594 18634 3654
rect 18520 3554 18556 3594
rect 18596 3554 18634 3594
rect 18520 3494 18634 3554
rect 18520 3454 18556 3494
rect 18596 3454 18634 3494
rect 18520 3384 18634 3454
rect 18664 3794 18778 3864
rect 18664 3754 18700 3794
rect 18740 3754 18778 3794
rect 18664 3694 18778 3754
rect 18664 3654 18700 3694
rect 18740 3654 18778 3694
rect 18664 3594 18778 3654
rect 18664 3554 18700 3594
rect 18740 3554 18778 3594
rect 18664 3494 18778 3554
rect 18664 3454 18700 3494
rect 18740 3454 18778 3494
rect 18664 3384 18778 3454
rect 18808 3794 18922 3864
rect 18808 3754 18844 3794
rect 18884 3754 18922 3794
rect 18808 3694 18922 3754
rect 18808 3654 18844 3694
rect 18884 3654 18922 3694
rect 18808 3594 18922 3654
rect 18808 3554 18844 3594
rect 18884 3554 18922 3594
rect 18808 3494 18922 3554
rect 18808 3454 18844 3494
rect 18884 3454 18922 3494
rect 18808 3384 18922 3454
rect 18952 3794 19066 3864
rect 18952 3754 18988 3794
rect 19028 3754 19066 3794
rect 18952 3694 19066 3754
rect 18952 3654 18988 3694
rect 19028 3654 19066 3694
rect 18952 3594 19066 3654
rect 18952 3554 18988 3594
rect 19028 3554 19066 3594
rect 18952 3494 19066 3554
rect 18952 3454 18988 3494
rect 19028 3454 19066 3494
rect 18952 3384 19066 3454
rect 19096 3794 19210 3864
rect 19096 3754 19132 3794
rect 19172 3754 19210 3794
rect 19096 3694 19210 3754
rect 19096 3654 19132 3694
rect 19172 3654 19210 3694
rect 19096 3594 19210 3654
rect 19096 3554 19132 3594
rect 19172 3554 19210 3594
rect 19096 3494 19210 3554
rect 19096 3454 19132 3494
rect 19172 3454 19210 3494
rect 19096 3384 19210 3454
rect 19240 3794 19354 3864
rect 19240 3754 19276 3794
rect 19316 3754 19354 3794
rect 19240 3694 19354 3754
rect 19240 3654 19276 3694
rect 19316 3654 19354 3694
rect 19240 3594 19354 3654
rect 19240 3554 19276 3594
rect 19316 3554 19354 3594
rect 19240 3494 19354 3554
rect 19240 3454 19276 3494
rect 19316 3454 19354 3494
rect 19240 3384 19354 3454
rect 19384 3794 19498 3864
rect 19384 3754 19420 3794
rect 19460 3754 19498 3794
rect 19384 3694 19498 3754
rect 19384 3654 19420 3694
rect 19460 3654 19498 3694
rect 19384 3594 19498 3654
rect 19384 3554 19420 3594
rect 19460 3554 19498 3594
rect 19384 3494 19498 3554
rect 19384 3454 19420 3494
rect 19460 3454 19498 3494
rect 19384 3384 19498 3454
rect 19528 3794 19642 3864
rect 19528 3754 19564 3794
rect 19604 3754 19642 3794
rect 19528 3694 19642 3754
rect 19528 3654 19564 3694
rect 19604 3654 19642 3694
rect 19528 3594 19642 3654
rect 19528 3554 19564 3594
rect 19604 3554 19642 3594
rect 19528 3494 19642 3554
rect 19528 3454 19564 3494
rect 19604 3454 19642 3494
rect 19528 3384 19642 3454
rect 19672 3794 19786 3864
rect 19672 3754 19708 3794
rect 19748 3754 19786 3794
rect 19672 3694 19786 3754
rect 19672 3654 19708 3694
rect 19748 3654 19786 3694
rect 19672 3594 19786 3654
rect 19672 3554 19708 3594
rect 19748 3554 19786 3594
rect 19672 3494 19786 3554
rect 19672 3454 19708 3494
rect 19748 3454 19786 3494
rect 19672 3384 19786 3454
rect 19816 3794 19930 3864
rect 19816 3754 19852 3794
rect 19892 3754 19930 3794
rect 19816 3694 19930 3754
rect 19816 3654 19852 3694
rect 19892 3654 19930 3694
rect 19816 3594 19930 3654
rect 19816 3554 19852 3594
rect 19892 3554 19930 3594
rect 19816 3494 19930 3554
rect 19816 3454 19852 3494
rect 19892 3454 19930 3494
rect 19816 3384 19930 3454
rect 19960 3794 20072 3864
rect 19960 3754 19996 3794
rect 20036 3754 20072 3794
rect 19960 3694 20072 3754
rect 19960 3654 19996 3694
rect 20036 3654 20072 3694
rect 19960 3594 20072 3654
rect 19960 3554 19996 3594
rect 20036 3554 20072 3594
rect 19960 3494 20072 3554
rect 19960 3454 19996 3494
rect 20036 3454 20072 3494
rect 19960 3384 20072 3454
rect 664 578 776 648
rect 664 538 700 578
rect 740 538 776 578
rect 664 478 776 538
rect 664 438 700 478
rect 740 438 776 478
rect 664 378 776 438
rect 664 338 700 378
rect 740 338 776 378
rect 664 278 776 338
rect 664 238 700 278
rect 740 238 776 278
rect 664 168 776 238
rect 806 578 920 648
rect 806 538 844 578
rect 884 538 920 578
rect 806 478 920 538
rect 806 438 844 478
rect 884 438 920 478
rect 806 378 920 438
rect 806 338 844 378
rect 884 338 920 378
rect 806 278 920 338
rect 806 238 844 278
rect 884 238 920 278
rect 806 168 920 238
rect 950 578 1064 648
rect 950 538 988 578
rect 1028 538 1064 578
rect 950 478 1064 538
rect 950 438 988 478
rect 1028 438 1064 478
rect 950 378 1064 438
rect 950 338 988 378
rect 1028 338 1064 378
rect 950 278 1064 338
rect 950 238 988 278
rect 1028 238 1064 278
rect 950 168 1064 238
rect 1240 578 1352 648
rect 1240 538 1276 578
rect 1316 538 1352 578
rect 1240 478 1352 538
rect 1240 438 1276 478
rect 1316 438 1352 478
rect 1240 378 1352 438
rect 1240 338 1276 378
rect 1316 338 1352 378
rect 1240 278 1352 338
rect 1240 238 1276 278
rect 1316 238 1352 278
rect 1240 168 1352 238
rect 1382 578 1496 648
rect 1382 538 1420 578
rect 1460 538 1496 578
rect 1382 478 1496 538
rect 1382 438 1420 478
rect 1460 438 1496 478
rect 1382 378 1496 438
rect 1382 338 1420 378
rect 1460 338 1496 378
rect 1382 278 1496 338
rect 1382 238 1420 278
rect 1460 238 1496 278
rect 1382 168 1496 238
rect 1526 578 1640 648
rect 1526 538 1564 578
rect 1604 538 1640 578
rect 1526 478 1640 538
rect 1526 438 1564 478
rect 1604 438 1640 478
rect 1526 378 1640 438
rect 1526 338 1564 378
rect 1604 338 1640 378
rect 1526 278 1640 338
rect 1526 238 1564 278
rect 1604 238 1640 278
rect 1526 168 1640 238
rect 1816 578 1928 648
rect 1816 538 1852 578
rect 1892 538 1928 578
rect 1816 478 1928 538
rect 1816 438 1852 478
rect 1892 438 1928 478
rect 1816 378 1928 438
rect 1816 338 1852 378
rect 1892 338 1928 378
rect 1816 278 1928 338
rect 1816 238 1852 278
rect 1892 238 1928 278
rect 1816 168 1928 238
rect 1958 578 2072 648
rect 1958 538 1996 578
rect 2036 538 2072 578
rect 1958 478 2072 538
rect 1958 438 1996 478
rect 2036 438 2072 478
rect 1958 378 2072 438
rect 1958 338 1996 378
rect 2036 338 2072 378
rect 1958 278 2072 338
rect 1958 238 1996 278
rect 2036 238 2072 278
rect 1958 168 2072 238
rect 2102 578 2216 648
rect 2102 538 2140 578
rect 2180 538 2216 578
rect 2102 478 2216 538
rect 2102 438 2140 478
rect 2180 438 2216 478
rect 2102 378 2216 438
rect 2102 338 2140 378
rect 2180 338 2216 378
rect 2102 278 2216 338
rect 2102 238 2140 278
rect 2180 238 2216 278
rect 2102 168 2216 238
rect 2968 578 3080 648
rect 2968 538 3004 578
rect 3044 538 3080 578
rect 2968 478 3080 538
rect 2968 438 3004 478
rect 3044 438 3080 478
rect 2968 378 3080 438
rect 2968 338 3004 378
rect 3044 338 3080 378
rect 2968 278 3080 338
rect 2968 238 3004 278
rect 3044 238 3080 278
rect 2968 168 3080 238
rect 3110 578 3224 648
rect 3110 538 3148 578
rect 3188 538 3224 578
rect 3110 478 3224 538
rect 3110 438 3148 478
rect 3188 438 3224 478
rect 3110 378 3224 438
rect 3110 338 3148 378
rect 3188 338 3224 378
rect 3110 278 3224 338
rect 3110 238 3148 278
rect 3188 238 3224 278
rect 3110 168 3224 238
rect 3254 578 3368 648
rect 3254 538 3292 578
rect 3332 538 3368 578
rect 3254 478 3368 538
rect 3254 438 3292 478
rect 3332 438 3368 478
rect 3254 378 3368 438
rect 3254 338 3292 378
rect 3332 338 3368 378
rect 3254 278 3368 338
rect 3254 238 3292 278
rect 3332 238 3368 278
rect 3254 168 3368 238
rect 3544 578 3656 648
rect 3544 538 3580 578
rect 3620 538 3656 578
rect 3544 478 3656 538
rect 3544 438 3580 478
rect 3620 438 3656 478
rect 3544 378 3656 438
rect 3544 338 3580 378
rect 3620 338 3656 378
rect 3544 278 3656 338
rect 3544 238 3580 278
rect 3620 238 3656 278
rect 3544 168 3656 238
rect 3686 578 3800 648
rect 3686 538 3724 578
rect 3764 538 3800 578
rect 3686 478 3800 538
rect 3686 438 3724 478
rect 3764 438 3800 478
rect 3686 378 3800 438
rect 3686 338 3724 378
rect 3764 338 3800 378
rect 3686 278 3800 338
rect 3686 238 3724 278
rect 3764 238 3800 278
rect 3686 168 3800 238
rect 3830 578 3944 648
rect 3830 538 3868 578
rect 3908 538 3944 578
rect 3830 478 3944 538
rect 3830 438 3868 478
rect 3908 438 3944 478
rect 3830 378 3944 438
rect 3830 338 3868 378
rect 3908 338 3944 378
rect 3830 278 3944 338
rect 3830 238 3868 278
rect 3908 238 3944 278
rect 3830 168 3944 238
rect 4120 578 4232 648
rect 4120 538 4156 578
rect 4196 538 4232 578
rect 4120 478 4232 538
rect 4120 438 4156 478
rect 4196 438 4232 478
rect 4120 378 4232 438
rect 4120 338 4156 378
rect 4196 338 4232 378
rect 4120 278 4232 338
rect 4120 238 4156 278
rect 4196 238 4232 278
rect 4120 168 4232 238
rect 4262 578 4376 648
rect 4262 538 4300 578
rect 4340 538 4376 578
rect 4262 478 4376 538
rect 4262 438 4300 478
rect 4340 438 4376 478
rect 4262 378 4376 438
rect 4262 338 4300 378
rect 4340 338 4376 378
rect 4262 278 4376 338
rect 4262 238 4300 278
rect 4340 238 4376 278
rect 4262 168 4376 238
rect 4406 578 4520 648
rect 4406 538 4444 578
rect 4484 538 4520 578
rect 4406 478 4520 538
rect 5848 578 5960 648
rect 5848 538 5884 578
rect 5924 538 5960 578
rect 4406 438 4444 478
rect 4484 438 4520 478
rect 4406 378 4520 438
rect 4406 338 4444 378
rect 4484 338 4520 378
rect 4406 278 4520 338
rect 5848 478 5960 538
rect 5848 438 5884 478
rect 5924 438 5960 478
rect 5848 378 5960 438
rect 5848 338 5884 378
rect 5924 338 5960 378
rect 4406 238 4444 278
rect 4484 238 4520 278
rect 4406 168 4520 238
rect 5848 278 5960 338
rect 5848 238 5884 278
rect 5924 238 5960 278
rect 5848 168 5960 238
rect 5990 578 6104 648
rect 5990 538 6028 578
rect 6068 538 6104 578
rect 5990 478 6104 538
rect 5990 438 6028 478
rect 6068 438 6104 478
rect 5990 378 6104 438
rect 5990 338 6028 378
rect 6068 338 6104 378
rect 5990 278 6104 338
rect 5990 238 6028 278
rect 6068 238 6104 278
rect 5990 168 6104 238
rect 6134 578 6248 648
rect 6134 538 6172 578
rect 6212 538 6248 578
rect 6134 478 6248 538
rect 6134 438 6172 478
rect 6212 438 6248 478
rect 6134 378 6248 438
rect 6134 338 6172 378
rect 6212 338 6248 378
rect 6134 278 6248 338
rect 6134 238 6172 278
rect 6212 238 6248 278
rect 6134 168 6248 238
rect 6424 578 6536 648
rect 6424 538 6460 578
rect 6500 538 6536 578
rect 6424 478 6536 538
rect 6424 438 6460 478
rect 6500 438 6536 478
rect 6424 378 6536 438
rect 6424 338 6460 378
rect 6500 338 6536 378
rect 6424 278 6536 338
rect 6424 238 6460 278
rect 6500 238 6536 278
rect 6424 168 6536 238
rect 6566 578 6680 648
rect 6566 538 6604 578
rect 6644 538 6680 578
rect 6566 478 6680 538
rect 6566 438 6604 478
rect 6644 438 6680 478
rect 6566 378 6680 438
rect 6566 338 6604 378
rect 6644 338 6680 378
rect 6566 278 6680 338
rect 6566 238 6604 278
rect 6644 238 6680 278
rect 6566 168 6680 238
rect 6710 578 6824 648
rect 6710 538 6748 578
rect 6788 538 6824 578
rect 6710 478 6824 538
rect 6710 438 6748 478
rect 6788 438 6824 478
rect 6710 378 6824 438
rect 6710 338 6748 378
rect 6788 338 6824 378
rect 6710 278 6824 338
rect 6710 238 6748 278
rect 6788 238 6824 278
rect 6710 168 6824 238
rect 7000 578 7112 648
rect 7000 538 7036 578
rect 7076 538 7112 578
rect 7000 478 7112 538
rect 7000 438 7036 478
rect 7076 438 7112 478
rect 7000 378 7112 438
rect 7000 338 7036 378
rect 7076 338 7112 378
rect 7000 278 7112 338
rect 7000 238 7036 278
rect 7076 238 7112 278
rect 7000 168 7112 238
rect 7142 578 7256 648
rect 7142 538 7180 578
rect 7220 538 7256 578
rect 7142 478 7256 538
rect 7142 438 7180 478
rect 7220 438 7256 478
rect 7142 378 7256 438
rect 7142 338 7180 378
rect 7220 338 7256 378
rect 7142 278 7256 338
rect 7142 238 7180 278
rect 7220 238 7256 278
rect 7142 168 7256 238
rect 7286 578 7400 648
rect 7286 538 7324 578
rect 7364 538 7400 578
rect 7286 478 7400 538
rect 7286 438 7324 478
rect 7364 438 7400 478
rect 7286 378 7400 438
rect 7286 338 7324 378
rect 7364 338 7400 378
rect 7286 278 7400 338
rect 7286 238 7324 278
rect 7364 238 7400 278
rect 7286 168 7400 238
rect 7576 578 7688 648
rect 7576 538 7612 578
rect 7652 538 7688 578
rect 7576 478 7688 538
rect 7576 438 7612 478
rect 7652 438 7688 478
rect 7576 378 7688 438
rect 7576 338 7612 378
rect 7652 338 7688 378
rect 7576 278 7688 338
rect 7576 238 7612 278
rect 7652 238 7688 278
rect 7576 168 7688 238
rect 7718 578 7832 648
rect 7718 538 7756 578
rect 7796 538 7832 578
rect 7718 478 7832 538
rect 7718 438 7756 478
rect 7796 438 7832 478
rect 7718 378 7832 438
rect 7718 338 7756 378
rect 7796 338 7832 378
rect 7718 278 7832 338
rect 7718 238 7756 278
rect 7796 238 7832 278
rect 7718 168 7832 238
rect 7862 578 7976 648
rect 7862 538 7900 578
rect 7940 538 7976 578
rect 7862 478 7976 538
rect 7862 438 7900 478
rect 7940 438 7976 478
rect 7862 378 7976 438
rect 7862 338 7900 378
rect 7940 338 7976 378
rect 7862 278 7976 338
rect 7862 238 7900 278
rect 7940 238 7976 278
rect 7862 168 7976 238
rect 8152 578 8264 648
rect 8152 538 8188 578
rect 8228 538 8264 578
rect 8152 478 8264 538
rect 8152 438 8188 478
rect 8228 438 8264 478
rect 8152 378 8264 438
rect 8152 338 8188 378
rect 8228 338 8264 378
rect 8152 278 8264 338
rect 8152 238 8188 278
rect 8228 238 8264 278
rect 8152 168 8264 238
rect 8294 578 8408 648
rect 8294 538 8332 578
rect 8372 538 8408 578
rect 8294 478 8408 538
rect 8294 438 8332 478
rect 8372 438 8408 478
rect 8294 378 8408 438
rect 8294 338 8332 378
rect 8372 338 8408 378
rect 8294 278 8408 338
rect 8294 238 8332 278
rect 8372 238 8408 278
rect 8294 168 8408 238
rect 8438 578 8552 648
rect 8438 538 8476 578
rect 8516 538 8552 578
rect 8438 478 8552 538
rect 9304 578 9416 648
rect 9304 538 9340 578
rect 9380 538 9416 578
rect 8438 438 8476 478
rect 8516 438 8552 478
rect 8438 378 8552 438
rect 8438 338 8476 378
rect 8516 338 8552 378
rect 8438 278 8552 338
rect 9304 478 9416 538
rect 9304 438 9340 478
rect 9380 438 9416 478
rect 9304 378 9416 438
rect 9304 338 9340 378
rect 9380 338 9416 378
rect 8438 238 8476 278
rect 8516 238 8552 278
rect 8438 168 8552 238
rect 9304 278 9416 338
rect 9304 238 9340 278
rect 9380 238 9416 278
rect 9304 168 9416 238
rect 9446 578 9560 648
rect 9446 538 9484 578
rect 9524 538 9560 578
rect 9446 478 9560 538
rect 9446 438 9484 478
rect 9524 438 9560 478
rect 9446 378 9560 438
rect 9446 338 9484 378
rect 9524 338 9560 378
rect 9446 278 9560 338
rect 9446 238 9484 278
rect 9524 238 9560 278
rect 9446 168 9560 238
rect 9590 578 9704 648
rect 9590 538 9628 578
rect 9668 538 9704 578
rect 9590 478 9704 538
rect 9590 438 9628 478
rect 9668 438 9704 478
rect 9590 378 9704 438
rect 9590 338 9628 378
rect 9668 338 9704 378
rect 9590 278 9704 338
rect 9590 238 9628 278
rect 9668 238 9704 278
rect 9590 168 9704 238
rect 9880 578 9992 648
rect 9880 538 9916 578
rect 9956 538 9992 578
rect 9880 478 9992 538
rect 9880 438 9916 478
rect 9956 438 9992 478
rect 9880 378 9992 438
rect 9880 338 9916 378
rect 9956 338 9992 378
rect 9880 278 9992 338
rect 9880 238 9916 278
rect 9956 238 9992 278
rect 9880 168 9992 238
rect 10022 578 10136 648
rect 10022 538 10060 578
rect 10100 538 10136 578
rect 10022 478 10136 538
rect 10022 438 10060 478
rect 10100 438 10136 478
rect 10022 378 10136 438
rect 10022 338 10060 378
rect 10100 338 10136 378
rect 10022 278 10136 338
rect 10022 238 10060 278
rect 10100 238 10136 278
rect 10022 168 10136 238
rect 10166 578 10280 648
rect 10166 538 10204 578
rect 10244 538 10280 578
rect 10166 478 10280 538
rect 10166 438 10204 478
rect 10244 438 10280 478
rect 10166 378 10280 438
rect 10166 338 10204 378
rect 10244 338 10280 378
rect 10166 278 10280 338
rect 10166 238 10204 278
rect 10244 238 10280 278
rect 10166 168 10280 238
rect 10456 578 10568 648
rect 10456 538 10492 578
rect 10532 538 10568 578
rect 10456 478 10568 538
rect 10456 438 10492 478
rect 10532 438 10568 478
rect 10456 378 10568 438
rect 10456 338 10492 378
rect 10532 338 10568 378
rect 10456 278 10568 338
rect 10456 238 10492 278
rect 10532 238 10568 278
rect 10456 168 10568 238
rect 10598 578 10712 648
rect 10598 538 10636 578
rect 10676 538 10712 578
rect 10598 478 10712 538
rect 10598 438 10636 478
rect 10676 438 10712 478
rect 10598 378 10712 438
rect 10598 338 10636 378
rect 10676 338 10712 378
rect 10598 278 10712 338
rect 10598 238 10636 278
rect 10676 238 10712 278
rect 10598 168 10712 238
rect 10742 578 10856 648
rect 10742 538 10780 578
rect 10820 538 10856 578
rect 10742 478 10856 538
rect 10742 438 10780 478
rect 10820 438 10856 478
rect 10742 378 10856 438
rect 10742 338 10780 378
rect 10820 338 10856 378
rect 10742 278 10856 338
rect 10742 238 10780 278
rect 10820 238 10856 278
rect 10742 168 10856 238
rect 11032 578 11144 648
rect 11032 538 11068 578
rect 11108 538 11144 578
rect 11032 478 11144 538
rect 11032 438 11068 478
rect 11108 438 11144 478
rect 11032 378 11144 438
rect 11032 338 11068 378
rect 11108 338 11144 378
rect 11032 278 11144 338
rect 11032 238 11068 278
rect 11108 238 11144 278
rect 11032 168 11144 238
rect 11174 578 11288 648
rect 11174 538 11212 578
rect 11252 538 11288 578
rect 11174 478 11288 538
rect 11174 438 11212 478
rect 11252 438 11288 478
rect 11174 378 11288 438
rect 11174 338 11212 378
rect 11252 338 11288 378
rect 11174 278 11288 338
rect 11174 238 11212 278
rect 11252 238 11288 278
rect 11174 168 11288 238
rect 11318 578 11432 648
rect 11318 538 11356 578
rect 11396 538 11432 578
rect 11318 478 11432 538
rect 11318 438 11356 478
rect 11396 438 11432 478
rect 11318 378 11432 438
rect 11318 338 11356 378
rect 11396 338 11432 378
rect 11318 278 11432 338
rect 11318 238 11356 278
rect 11396 238 11432 278
rect 11318 168 11432 238
rect 11896 578 12008 648
rect 11896 538 11932 578
rect 11972 538 12008 578
rect 11896 478 12008 538
rect 11896 438 11932 478
rect 11972 438 12008 478
rect 11896 378 12008 438
rect 11896 338 11932 378
rect 11972 338 12008 378
rect 11896 278 12008 338
rect 11896 238 11932 278
rect 11972 238 12008 278
rect 11896 168 12008 238
rect 12038 578 12152 648
rect 12038 538 12076 578
rect 12116 538 12152 578
rect 12038 478 12152 538
rect 12038 438 12076 478
rect 12116 438 12152 478
rect 12038 378 12152 438
rect 12038 338 12076 378
rect 12116 338 12152 378
rect 12038 278 12152 338
rect 12038 238 12076 278
rect 12116 238 12152 278
rect 12038 168 12152 238
rect 12182 578 12296 648
rect 12182 538 12220 578
rect 12260 538 12296 578
rect 12182 478 12296 538
rect 12182 438 12220 478
rect 12260 438 12296 478
rect 12182 378 12296 438
rect 12182 338 12220 378
rect 12260 338 12296 378
rect 12182 278 12296 338
rect 12182 238 12220 278
rect 12260 238 12296 278
rect 12182 168 12296 238
rect 12472 578 12584 648
rect 12472 538 12508 578
rect 12548 538 12584 578
rect 12472 478 12584 538
rect 12472 438 12508 478
rect 12548 438 12584 478
rect 12472 378 12584 438
rect 12472 338 12508 378
rect 12548 338 12584 378
rect 12472 278 12584 338
rect 12472 238 12508 278
rect 12548 238 12584 278
rect 12472 168 12584 238
rect 12614 578 12728 648
rect 12614 538 12652 578
rect 12692 538 12728 578
rect 12614 478 12728 538
rect 12614 438 12652 478
rect 12692 438 12728 478
rect 12614 378 12728 438
rect 12614 338 12652 378
rect 12692 338 12728 378
rect 12614 278 12728 338
rect 12614 238 12652 278
rect 12692 238 12728 278
rect 12614 168 12728 238
rect 12758 578 12872 648
rect 12758 538 12796 578
rect 12836 538 12872 578
rect 12758 478 12872 538
rect 12758 438 12796 478
rect 12836 438 12872 478
rect 12758 378 12872 438
rect 12758 338 12796 378
rect 12836 338 12872 378
rect 12758 278 12872 338
rect 12758 238 12796 278
rect 12836 238 12872 278
rect 12758 168 12872 238
rect 13048 578 13160 648
rect 13048 538 13084 578
rect 13124 538 13160 578
rect 13048 478 13160 538
rect 13048 438 13084 478
rect 13124 438 13160 478
rect 13048 378 13160 438
rect 13048 338 13084 378
rect 13124 338 13160 378
rect 13048 278 13160 338
rect 13048 238 13084 278
rect 13124 238 13160 278
rect 13048 168 13160 238
rect 13190 578 13304 648
rect 13190 538 13228 578
rect 13268 538 13304 578
rect 13190 478 13304 538
rect 13190 438 13228 478
rect 13268 438 13304 478
rect 13190 378 13304 438
rect 13190 338 13228 378
rect 13268 338 13304 378
rect 13190 278 13304 338
rect 13190 238 13228 278
rect 13268 238 13304 278
rect 13190 168 13304 238
rect 13334 578 13448 648
rect 13334 538 13372 578
rect 13412 538 13448 578
rect 13334 478 13448 538
rect 13334 438 13372 478
rect 13412 438 13448 478
rect 13334 378 13448 438
rect 13334 338 13372 378
rect 13412 338 13448 378
rect 13334 278 13448 338
rect 13334 238 13372 278
rect 13412 238 13448 278
rect 13334 168 13448 238
rect 13624 578 13736 648
rect 13624 538 13660 578
rect 13700 538 13736 578
rect 13624 478 13736 538
rect 13624 438 13660 478
rect 13700 438 13736 478
rect 13624 378 13736 438
rect 13624 338 13660 378
rect 13700 338 13736 378
rect 13624 278 13736 338
rect 13624 238 13660 278
rect 13700 238 13736 278
rect 13624 168 13736 238
rect 13766 578 13880 648
rect 13766 538 13804 578
rect 13844 538 13880 578
rect 13766 478 13880 538
rect 13766 438 13804 478
rect 13844 438 13880 478
rect 13766 378 13880 438
rect 13766 338 13804 378
rect 13844 338 13880 378
rect 13766 278 13880 338
rect 13766 238 13804 278
rect 13844 238 13880 278
rect 13766 168 13880 238
rect 13910 578 14024 648
rect 13910 538 13948 578
rect 13988 538 14024 578
rect 13910 478 14024 538
rect 14776 578 14888 648
rect 14776 538 14812 578
rect 14852 538 14888 578
rect 13910 438 13948 478
rect 13988 438 14024 478
rect 13910 378 14024 438
rect 13910 338 13948 378
rect 13988 338 14024 378
rect 13910 278 14024 338
rect 14776 478 14888 538
rect 14776 438 14812 478
rect 14852 438 14888 478
rect 14776 378 14888 438
rect 14776 338 14812 378
rect 14852 338 14888 378
rect 13910 238 13948 278
rect 13988 238 14024 278
rect 13910 168 14024 238
rect 14776 278 14888 338
rect 14776 238 14812 278
rect 14852 238 14888 278
rect 14776 168 14888 238
rect 14918 578 15032 648
rect 14918 538 14956 578
rect 14996 538 15032 578
rect 14918 478 15032 538
rect 14918 438 14956 478
rect 14996 438 15032 478
rect 14918 378 15032 438
rect 14918 338 14956 378
rect 14996 338 15032 378
rect 14918 278 15032 338
rect 14918 238 14956 278
rect 14996 238 15032 278
rect 14918 168 15032 238
rect 15062 578 15176 648
rect 15062 538 15100 578
rect 15140 538 15176 578
rect 15062 478 15176 538
rect 15062 438 15100 478
rect 15140 438 15176 478
rect 15062 378 15176 438
rect 15062 338 15100 378
rect 15140 338 15176 378
rect 15062 278 15176 338
rect 15062 238 15100 278
rect 15140 238 15176 278
rect 15062 168 15176 238
rect 15352 578 15466 648
rect 15352 538 15388 578
rect 15428 538 15466 578
rect 15352 478 15466 538
rect 15352 438 15388 478
rect 15428 438 15466 478
rect 15352 378 15466 438
rect 15352 338 15388 378
rect 15428 338 15466 378
rect 15352 278 15466 338
rect 15352 238 15388 278
rect 15428 238 15466 278
rect 15352 168 15466 238
rect 15496 578 15610 648
rect 15496 538 15532 578
rect 15572 538 15610 578
rect 15496 478 15610 538
rect 15496 438 15532 478
rect 15572 438 15610 478
rect 15496 378 15610 438
rect 15496 338 15532 378
rect 15572 338 15610 378
rect 15496 278 15610 338
rect 15496 238 15532 278
rect 15572 238 15610 278
rect 15496 168 15610 238
rect 15640 578 15752 648
rect 15640 538 15676 578
rect 15716 538 15752 578
rect 15640 478 15752 538
rect 15640 438 15676 478
rect 15716 438 15752 478
rect 15640 378 15752 438
rect 15640 338 15676 378
rect 15716 338 15752 378
rect 15640 278 15752 338
rect 15640 238 15676 278
rect 15716 238 15752 278
rect 15640 168 15752 238
rect 15928 578 16040 648
rect 15928 538 15964 578
rect 16004 538 16040 578
rect 15928 478 16040 538
rect 15928 438 15964 478
rect 16004 438 16040 478
rect 15928 378 16040 438
rect 15928 338 15964 378
rect 16004 338 16040 378
rect 15928 278 16040 338
rect 15928 238 15964 278
rect 16004 238 16040 278
rect 15928 168 16040 238
rect 16070 578 16184 648
rect 16070 538 16108 578
rect 16148 538 16184 578
rect 16070 478 16184 538
rect 16070 438 16108 478
rect 16148 438 16184 478
rect 16070 378 16184 438
rect 16070 338 16108 378
rect 16148 338 16184 378
rect 16070 278 16184 338
rect 16070 238 16108 278
rect 16148 238 16184 278
rect 16070 168 16184 238
rect 16214 578 16328 648
rect 16214 538 16252 578
rect 16292 538 16328 578
rect 16214 478 16328 538
rect 16214 438 16252 478
rect 16292 438 16328 478
rect 16214 378 16328 438
rect 16214 338 16252 378
rect 16292 338 16328 378
rect 16214 278 16328 338
rect 16214 238 16252 278
rect 16292 238 16328 278
rect 16214 168 16328 238
rect 16358 578 16472 648
rect 16358 538 16396 578
rect 16436 538 16472 578
rect 16358 478 16472 538
rect 16358 438 16396 478
rect 16436 438 16472 478
rect 16358 378 16472 438
rect 16358 338 16396 378
rect 16436 338 16472 378
rect 16358 278 16472 338
rect 16358 238 16396 278
rect 16436 238 16472 278
rect 16358 168 16472 238
rect 16502 578 16616 648
rect 16502 538 16540 578
rect 16580 538 16616 578
rect 16502 478 16616 538
rect 17368 578 17480 648
rect 17368 538 17404 578
rect 17444 538 17480 578
rect 16502 438 16540 478
rect 16580 438 16616 478
rect 16502 378 16616 438
rect 16502 338 16540 378
rect 16580 338 16616 378
rect 16502 278 16616 338
rect 17368 478 17480 538
rect 17368 438 17404 478
rect 17444 438 17480 478
rect 17368 378 17480 438
rect 17368 338 17404 378
rect 17444 338 17480 378
rect 16502 238 16540 278
rect 16580 238 16616 278
rect 16502 168 16616 238
rect 17368 278 17480 338
rect 17368 238 17404 278
rect 17444 238 17480 278
rect 17368 168 17480 238
rect 17510 578 17624 648
rect 17510 538 17548 578
rect 17588 538 17624 578
rect 17510 478 17624 538
rect 17510 438 17548 478
rect 17588 438 17624 478
rect 17510 378 17624 438
rect 17510 338 17548 378
rect 17588 338 17624 378
rect 17510 278 17624 338
rect 17510 238 17548 278
rect 17588 238 17624 278
rect 17510 168 17624 238
rect 17654 578 17768 648
rect 17654 538 17692 578
rect 17732 538 17768 578
rect 17654 478 17768 538
rect 17654 438 17692 478
rect 17732 438 17768 478
rect 17654 378 17768 438
rect 17654 338 17692 378
rect 17732 338 17768 378
rect 17654 278 17768 338
rect 17654 238 17692 278
rect 17732 238 17768 278
rect 17654 168 17768 238
rect 17798 578 17912 648
rect 17798 538 17836 578
rect 17876 538 17912 578
rect 17798 478 17912 538
rect 17798 438 17836 478
rect 17876 438 17912 478
rect 17798 378 17912 438
rect 17798 338 17836 378
rect 17876 338 17912 378
rect 17798 278 17912 338
rect 17798 238 17836 278
rect 17876 238 17912 278
rect 17798 168 17912 238
rect 17942 578 18056 648
rect 17942 538 17980 578
rect 18020 538 18056 578
rect 17942 478 18056 538
rect 17942 438 17980 478
rect 18020 438 18056 478
rect 17942 378 18056 438
rect 17942 338 17980 378
rect 18020 338 18056 378
rect 17942 278 18056 338
rect 17942 238 17980 278
rect 18020 238 18056 278
rect 17942 168 18056 238
rect 18086 578 18200 648
rect 18086 538 18124 578
rect 18164 538 18200 578
rect 18086 478 18200 538
rect 18086 438 18124 478
rect 18164 438 18200 478
rect 18086 378 18200 438
rect 18086 338 18124 378
rect 18164 338 18200 378
rect 18086 278 18200 338
rect 18086 238 18124 278
rect 18164 238 18200 278
rect 18086 168 18200 238
rect 18230 578 18344 648
rect 18230 538 18268 578
rect 18308 538 18344 578
rect 18230 478 18344 538
rect 18230 438 18268 478
rect 18308 438 18344 478
rect 18230 378 18344 438
rect 18230 338 18268 378
rect 18308 338 18344 378
rect 18230 278 18344 338
rect 18230 238 18268 278
rect 18308 238 18344 278
rect 18230 168 18344 238
rect 18374 578 18488 648
rect 18374 538 18412 578
rect 18452 538 18488 578
rect 18374 478 18488 538
rect 18374 438 18412 478
rect 18452 438 18488 478
rect 18374 378 18488 438
rect 18374 338 18412 378
rect 18452 338 18488 378
rect 18374 278 18488 338
rect 18374 238 18412 278
rect 18452 238 18488 278
rect 18374 168 18488 238
rect 18518 578 18632 648
rect 18518 538 18556 578
rect 18596 538 18632 578
rect 18518 478 18632 538
rect 18518 438 18556 478
rect 18596 438 18632 478
rect 18518 378 18632 438
rect 18518 338 18556 378
rect 18596 338 18632 378
rect 18518 278 18632 338
rect 18518 238 18556 278
rect 18596 238 18632 278
rect 18518 168 18632 238
rect 18662 578 18776 648
rect 18662 538 18700 578
rect 18740 538 18776 578
rect 18662 478 18776 538
rect 18662 438 18700 478
rect 18740 438 18776 478
rect 18662 378 18776 438
rect 18662 338 18700 378
rect 18740 338 18776 378
rect 18662 278 18776 338
rect 18662 238 18700 278
rect 18740 238 18776 278
rect 18662 168 18776 238
rect 18806 578 18920 648
rect 18806 538 18844 578
rect 18884 538 18920 578
rect 18806 478 18920 538
rect 18806 438 18844 478
rect 18884 438 18920 478
rect 18806 378 18920 438
rect 18806 338 18844 378
rect 18884 338 18920 378
rect 18806 278 18920 338
rect 18806 238 18844 278
rect 18884 238 18920 278
rect 18806 168 18920 238
rect 18950 578 19064 648
rect 18950 538 18988 578
rect 19028 538 19064 578
rect 18950 478 19064 538
rect 18950 438 18988 478
rect 19028 438 19064 478
rect 18950 378 19064 438
rect 18950 338 18988 378
rect 19028 338 19064 378
rect 18950 278 19064 338
rect 18950 238 18988 278
rect 19028 238 19064 278
rect 18950 168 19064 238
rect 19094 578 19208 648
rect 19094 538 19132 578
rect 19172 538 19208 578
rect 19094 478 19208 538
rect 19094 438 19132 478
rect 19172 438 19208 478
rect 19094 378 19208 438
rect 19094 338 19132 378
rect 19172 338 19208 378
rect 19094 278 19208 338
rect 19094 238 19132 278
rect 19172 238 19208 278
rect 19094 168 19208 238
rect 19238 578 19352 648
rect 19238 538 19276 578
rect 19316 538 19352 578
rect 19238 478 19352 538
rect 19238 438 19276 478
rect 19316 438 19352 478
rect 19238 378 19352 438
rect 19238 338 19276 378
rect 19316 338 19352 378
rect 19238 278 19352 338
rect 19238 238 19276 278
rect 19316 238 19352 278
rect 19238 168 19352 238
rect 19382 578 19496 648
rect 19382 538 19420 578
rect 19460 538 19496 578
rect 19382 478 19496 538
rect 19382 438 19420 478
rect 19460 438 19496 478
rect 19382 378 19496 438
rect 19382 338 19420 378
rect 19460 338 19496 378
rect 19382 278 19496 338
rect 19382 238 19420 278
rect 19460 238 19496 278
rect 19382 168 19496 238
rect 19526 578 19640 648
rect 19526 538 19564 578
rect 19604 538 19640 578
rect 19526 478 19640 538
rect 19526 438 19564 478
rect 19604 438 19640 478
rect 19526 378 19640 438
rect 19526 338 19564 378
rect 19604 338 19640 378
rect 19526 278 19640 338
rect 19526 238 19564 278
rect 19604 238 19640 278
rect 19526 168 19640 238
rect 19670 578 19784 648
rect 19670 538 19708 578
rect 19748 538 19784 578
rect 19670 478 19784 538
rect 19670 438 19708 478
rect 19748 438 19784 478
rect 19670 378 19784 438
rect 19670 338 19708 378
rect 19748 338 19784 378
rect 19670 278 19784 338
rect 19670 238 19708 278
rect 19748 238 19784 278
rect 19670 168 19784 238
rect 19814 578 19928 648
rect 19814 538 19852 578
rect 19892 538 19928 578
rect 19814 478 19928 538
rect 19814 438 19852 478
rect 19892 438 19928 478
rect 19814 378 19928 438
rect 19814 338 19852 378
rect 19892 338 19928 378
rect 19814 278 19928 338
rect 19814 238 19852 278
rect 19892 238 19928 278
rect 19814 168 19928 238
rect 19958 578 20072 648
rect 19958 538 19996 578
rect 20036 538 20072 578
rect 19958 478 20072 538
rect 19958 438 19996 478
rect 20036 438 20072 478
rect 19958 378 20072 438
rect 19958 338 19996 378
rect 20036 338 20072 378
rect 19958 278 20072 338
rect 19958 238 19996 278
rect 20036 238 20072 278
rect 19958 168 20072 238
rect 20102 578 20216 648
rect 20102 538 20140 578
rect 20180 538 20216 578
rect 20102 478 20216 538
rect 20102 438 20140 478
rect 20180 438 20216 478
rect 20102 378 20216 438
rect 20102 338 20140 378
rect 20180 338 20216 378
rect 20102 278 20216 338
rect 20102 238 20140 278
rect 20180 238 20216 278
rect 20102 168 20216 238
rect 20246 578 20360 648
rect 20246 538 20284 578
rect 20324 538 20360 578
rect 20246 478 20360 538
rect 20246 438 20284 478
rect 20324 438 20360 478
rect 20246 378 20360 438
rect 20246 338 20284 378
rect 20324 338 20360 378
rect 20246 278 20360 338
rect 20246 238 20284 278
rect 20324 238 20360 278
rect 20246 168 20360 238
rect 20390 578 20504 648
rect 20390 538 20428 578
rect 20468 538 20504 578
rect 20390 478 20504 538
rect 20390 438 20428 478
rect 20468 438 20504 478
rect 20390 378 20504 438
rect 20390 338 20428 378
rect 20468 338 20504 378
rect 20390 278 20504 338
rect 20390 238 20428 278
rect 20468 238 20504 278
rect 20390 168 20504 238
rect 20534 578 20648 648
rect 20534 538 20572 578
rect 20612 538 20648 578
rect 20534 478 20648 538
rect 20534 438 20572 478
rect 20612 438 20648 478
rect 20534 378 20648 438
rect 20534 338 20572 378
rect 20612 338 20648 378
rect 20534 278 20648 338
rect 20534 238 20572 278
rect 20612 238 20648 278
rect 20534 168 20648 238
rect 20678 578 20792 648
rect 20678 538 20716 578
rect 20756 538 20792 578
rect 20678 478 20792 538
rect 20678 438 20716 478
rect 20756 438 20792 478
rect 20678 378 20792 438
rect 20678 338 20716 378
rect 20756 338 20792 378
rect 20678 278 20792 338
rect 20678 238 20716 278
rect 20756 238 20792 278
rect 20678 168 20792 238
rect 20822 578 20936 648
rect 20822 538 20860 578
rect 20900 538 20936 578
rect 20822 478 20936 538
rect 20822 438 20860 478
rect 20900 438 20936 478
rect 20822 378 20936 438
rect 20822 338 20860 378
rect 20900 338 20936 378
rect 20822 278 20936 338
rect 20822 238 20860 278
rect 20900 238 20936 278
rect 20822 168 20936 238
<< ndiffc >>
rect 700 2574 740 2614
rect 700 2474 740 2514
rect 844 2574 884 2614
rect 844 2474 884 2514
rect 988 2574 1028 2614
rect 988 2474 1028 2514
rect 1276 2574 1316 2614
rect 1276 2474 1316 2514
rect 1420 2574 1460 2614
rect 1420 2474 1460 2514
rect 1564 2574 1604 2614
rect 1564 2474 1604 2514
rect 1852 2574 1892 2614
rect 1852 2474 1892 2514
rect 1996 2574 2036 2614
rect 1996 2474 2036 2514
rect 2140 2574 2180 2614
rect 2140 2474 2180 2514
rect 2428 2574 2468 2614
rect 2428 2474 2468 2514
rect 2572 2574 2612 2614
rect 2572 2474 2612 2514
rect 2716 2574 2756 2614
rect 2716 2474 2756 2514
rect 3004 2574 3044 2614
rect 3004 2474 3044 2514
rect 3148 2574 3188 2614
rect 3148 2474 3188 2514
rect 3292 2574 3332 2614
rect 3292 2474 3332 2514
rect 4156 2574 4196 2614
rect 4156 2474 4196 2514
rect 4300 2574 4340 2614
rect 4300 2474 4340 2514
rect 4444 2574 4484 2614
rect 4444 2474 4484 2514
rect 4732 2574 4772 2614
rect 4732 2474 4772 2514
rect 4876 2574 4916 2614
rect 4876 2474 4916 2514
rect 5020 2574 5060 2614
rect 5020 2474 5060 2514
rect 5308 2574 5348 2614
rect 5308 2474 5348 2514
rect 5452 2574 5492 2614
rect 5452 2474 5492 2514
rect 5596 2574 5636 2614
rect 5596 2474 5636 2514
rect 5884 2574 5924 2614
rect 5884 2474 5924 2514
rect 6028 2574 6068 2614
rect 6028 2474 6068 2514
rect 6172 2574 6212 2614
rect 6172 2474 6212 2514
rect 6460 2574 6500 2614
rect 6460 2474 6500 2514
rect 6604 2574 6644 2614
rect 6604 2474 6644 2514
rect 6748 2574 6788 2614
rect 6748 2474 6788 2514
rect 7612 2574 7652 2614
rect 7612 2474 7652 2514
rect 7756 2574 7796 2614
rect 7756 2474 7796 2514
rect 7900 2574 7940 2614
rect 7900 2474 7940 2514
rect 8188 2574 8228 2614
rect 8188 2474 8228 2514
rect 8332 2574 8372 2614
rect 8332 2474 8372 2514
rect 8476 2574 8516 2614
rect 8476 2474 8516 2514
rect 8764 2574 8804 2614
rect 8764 2474 8804 2514
rect 8908 2574 8948 2614
rect 8908 2474 8948 2514
rect 9052 2574 9092 2614
rect 9052 2474 9092 2514
rect 9340 2574 9380 2614
rect 9340 2474 9380 2514
rect 9484 2574 9524 2614
rect 9484 2474 9524 2514
rect 9628 2574 9668 2614
rect 9628 2474 9668 2514
rect 10204 2574 10244 2614
rect 10204 2474 10244 2514
rect 10348 2574 10388 2614
rect 10348 2474 10388 2514
rect 10492 2574 10532 2614
rect 10492 2474 10532 2514
rect 10780 2574 10820 2614
rect 10780 2474 10820 2514
rect 10924 2574 10964 2614
rect 10924 2474 10964 2514
rect 11068 2574 11108 2614
rect 11068 2474 11108 2514
rect 11932 2574 11972 2614
rect 11932 2474 11972 2514
rect 12076 2574 12116 2614
rect 12076 2474 12116 2514
rect 12220 2574 12260 2614
rect 12220 2474 12260 2514
rect 12508 2574 12548 2614
rect 12508 2474 12548 2514
rect 12652 2574 12692 2614
rect 12652 2474 12692 2514
rect 12796 2574 12836 2614
rect 12796 2474 12836 2514
rect 13660 2574 13700 2614
rect 13660 2474 13700 2514
rect 13804 2574 13844 2614
rect 13804 2474 13844 2514
rect 13948 2574 13988 2614
rect 13948 2474 13988 2514
rect 14236 2574 14276 2614
rect 14236 2474 14276 2514
rect 14380 2574 14420 2614
rect 14380 2474 14420 2514
rect 14524 2574 14564 2614
rect 14524 2474 14564 2514
rect 14812 2574 14852 2614
rect 14812 2474 14852 2514
rect 14956 2574 14996 2614
rect 14956 2474 14996 2514
rect 15100 2574 15140 2614
rect 15100 2474 15140 2514
rect 16540 2574 16580 2614
rect 16540 2474 16580 2514
rect 16684 2574 16724 2614
rect 16684 2474 16724 2514
rect 16828 2574 16868 2614
rect 16828 2474 16868 2514
rect 16972 2574 17012 2614
rect 16972 2474 17012 2514
rect 17116 2574 17156 2614
rect 17116 2474 17156 2514
rect 17260 2574 17300 2614
rect 17260 2474 17300 2514
rect 17404 2574 17444 2614
rect 17404 2474 17444 2514
rect 17548 2574 17588 2614
rect 17548 2474 17588 2514
rect 17692 2574 17732 2614
rect 17692 2474 17732 2514
rect 17836 2574 17876 2614
rect 17836 2474 17876 2514
rect 17980 2574 18020 2614
rect 17980 2474 18020 2514
rect 18124 2574 18164 2614
rect 18124 2474 18164 2514
rect 18268 2574 18308 2614
rect 18268 2474 18308 2514
rect 18412 2574 18452 2614
rect 18412 2474 18452 2514
rect 18556 2574 18596 2614
rect 18556 2474 18596 2514
rect 18700 2574 18740 2614
rect 18700 2474 18740 2514
rect 18844 2574 18884 2614
rect 18844 2474 18884 2514
rect 18988 2574 19028 2614
rect 18988 2474 19028 2514
rect 19132 2574 19172 2614
rect 19132 2474 19172 2514
rect 19276 2574 19316 2614
rect 19276 2474 19316 2514
rect 19420 2574 19460 2614
rect 19420 2474 19460 2514
rect 19564 2574 19604 2614
rect 19564 2474 19604 2514
rect 19708 2574 19748 2614
rect 19708 2474 19748 2514
rect 19852 2574 19892 2614
rect 19852 2474 19892 2514
rect 19996 2574 20036 2614
rect 19996 2474 20036 2514
rect 700 1518 740 1558
rect 700 1418 740 1458
rect 844 1518 884 1558
rect 844 1418 884 1458
rect 988 1518 1028 1558
rect 988 1418 1028 1458
rect 1276 1518 1316 1558
rect 1276 1418 1316 1458
rect 1420 1518 1460 1558
rect 1420 1418 1460 1458
rect 1564 1518 1604 1558
rect 1564 1418 1604 1458
rect 1852 1518 1892 1558
rect 1852 1418 1892 1458
rect 1996 1518 2036 1558
rect 1996 1418 2036 1458
rect 2140 1518 2180 1558
rect 2140 1418 2180 1458
rect 3004 1518 3044 1558
rect 3004 1418 3044 1458
rect 3148 1518 3188 1558
rect 3148 1418 3188 1458
rect 3292 1518 3332 1558
rect 3292 1418 3332 1458
rect 3580 1518 3620 1558
rect 3580 1418 3620 1458
rect 3724 1518 3764 1558
rect 3724 1418 3764 1458
rect 3868 1518 3908 1558
rect 3868 1418 3908 1458
rect 4156 1518 4196 1558
rect 4156 1418 4196 1458
rect 4300 1518 4340 1558
rect 4300 1418 4340 1458
rect 4444 1518 4484 1558
rect 4444 1418 4484 1458
rect 5884 1518 5924 1558
rect 5884 1418 5924 1458
rect 6028 1518 6068 1558
rect 6028 1418 6068 1458
rect 6172 1518 6212 1558
rect 6172 1418 6212 1458
rect 6460 1518 6500 1558
rect 6460 1418 6500 1458
rect 6604 1518 6644 1558
rect 6604 1418 6644 1458
rect 6748 1518 6788 1558
rect 6748 1418 6788 1458
rect 7036 1518 7076 1558
rect 7036 1418 7076 1458
rect 7180 1518 7220 1558
rect 7180 1418 7220 1458
rect 7324 1518 7364 1558
rect 7324 1418 7364 1458
rect 7612 1518 7652 1558
rect 7612 1418 7652 1458
rect 7756 1518 7796 1558
rect 7756 1418 7796 1458
rect 7900 1518 7940 1558
rect 7900 1418 7940 1458
rect 8188 1518 8228 1558
rect 8188 1418 8228 1458
rect 8332 1518 8372 1558
rect 8332 1418 8372 1458
rect 8476 1518 8516 1558
rect 8476 1418 8516 1458
rect 9340 1518 9380 1558
rect 9340 1418 9380 1458
rect 9484 1518 9524 1558
rect 9484 1418 9524 1458
rect 9628 1518 9668 1558
rect 9628 1418 9668 1458
rect 9916 1518 9956 1558
rect 9916 1418 9956 1458
rect 10060 1518 10100 1558
rect 10060 1418 10100 1458
rect 10204 1518 10244 1558
rect 10204 1418 10244 1458
rect 10492 1518 10532 1558
rect 10492 1418 10532 1458
rect 10636 1518 10676 1558
rect 10636 1418 10676 1458
rect 10780 1518 10820 1558
rect 10780 1418 10820 1458
rect 11068 1518 11108 1558
rect 11068 1418 11108 1458
rect 11212 1518 11252 1558
rect 11212 1418 11252 1458
rect 11356 1518 11396 1558
rect 11356 1418 11396 1458
rect 11932 1518 11972 1558
rect 11932 1418 11972 1458
rect 12076 1518 12116 1558
rect 12076 1418 12116 1458
rect 12220 1518 12260 1558
rect 12220 1418 12260 1458
rect 12508 1518 12548 1558
rect 12508 1418 12548 1458
rect 12652 1518 12692 1558
rect 12652 1418 12692 1458
rect 12796 1518 12836 1558
rect 12796 1418 12836 1458
rect 13084 1518 13124 1558
rect 13084 1418 13124 1458
rect 13228 1518 13268 1558
rect 13228 1418 13268 1458
rect 13372 1518 13412 1558
rect 13372 1418 13412 1458
rect 13660 1518 13700 1558
rect 13660 1418 13700 1458
rect 13804 1518 13844 1558
rect 13804 1418 13844 1458
rect 13948 1518 13988 1558
rect 13948 1418 13988 1458
rect 14812 1518 14852 1558
rect 14812 1418 14852 1458
rect 14956 1518 14996 1558
rect 14956 1418 14996 1458
rect 15100 1518 15140 1558
rect 15100 1418 15140 1458
rect 15388 1518 15428 1558
rect 15388 1418 15428 1458
rect 15532 1518 15572 1558
rect 15532 1418 15572 1458
rect 15676 1518 15716 1558
rect 15676 1418 15716 1458
rect 15964 1518 16004 1558
rect 15964 1418 16004 1458
rect 16108 1518 16148 1558
rect 16108 1418 16148 1458
rect 16252 1518 16292 1558
rect 16252 1418 16292 1458
rect 16396 1518 16436 1558
rect 16396 1418 16436 1458
rect 16540 1518 16580 1558
rect 16540 1418 16580 1458
rect 17404 1518 17444 1558
rect 17404 1418 17444 1458
rect 17548 1518 17588 1558
rect 17548 1418 17588 1458
rect 17692 1518 17732 1558
rect 17692 1418 17732 1458
rect 17836 1518 17876 1558
rect 17836 1418 17876 1458
rect 17980 1518 18020 1558
rect 17980 1418 18020 1458
rect 18124 1518 18164 1558
rect 18124 1418 18164 1458
rect 18268 1518 18308 1558
rect 18268 1418 18308 1458
rect 18412 1518 18452 1558
rect 18412 1418 18452 1458
rect 18556 1518 18596 1558
rect 18556 1418 18596 1458
rect 18700 1518 18740 1558
rect 18700 1418 18740 1458
rect 18844 1518 18884 1558
rect 18844 1418 18884 1458
rect 18988 1518 19028 1558
rect 18988 1418 19028 1458
rect 19132 1518 19172 1558
rect 19132 1418 19172 1458
rect 19276 1518 19316 1558
rect 19276 1418 19316 1458
rect 19420 1518 19460 1558
rect 19420 1418 19460 1458
rect 19564 1518 19604 1558
rect 19564 1418 19604 1458
rect 19708 1518 19748 1558
rect 19708 1418 19748 1458
rect 19852 1518 19892 1558
rect 19852 1418 19892 1458
rect 19996 1518 20036 1558
rect 19996 1418 20036 1458
rect 20140 1518 20180 1558
rect 20140 1418 20180 1458
rect 20284 1518 20324 1558
rect 20284 1418 20324 1458
rect 20428 1518 20468 1558
rect 20428 1418 20468 1458
rect 20572 1518 20612 1558
rect 20572 1418 20612 1458
rect 20716 1518 20756 1558
rect 20716 1418 20756 1458
rect 20860 1518 20900 1558
rect 20860 1418 20900 1458
<< pdiffc >>
rect 700 3754 740 3794
rect 700 3654 740 3694
rect 700 3554 740 3594
rect 700 3454 740 3494
rect 844 3754 884 3794
rect 844 3654 884 3694
rect 844 3554 884 3594
rect 844 3454 884 3494
rect 988 3754 1028 3794
rect 988 3654 1028 3694
rect 988 3554 1028 3594
rect 988 3454 1028 3494
rect 1276 3754 1316 3794
rect 1276 3654 1316 3694
rect 1276 3554 1316 3594
rect 1276 3454 1316 3494
rect 1420 3754 1460 3794
rect 1420 3654 1460 3694
rect 1420 3554 1460 3594
rect 1420 3454 1460 3494
rect 1564 3754 1604 3794
rect 1564 3654 1604 3694
rect 1564 3554 1604 3594
rect 1564 3454 1604 3494
rect 1852 3754 1892 3794
rect 1852 3654 1892 3694
rect 1852 3554 1892 3594
rect 1852 3454 1892 3494
rect 1996 3754 2036 3794
rect 1996 3654 2036 3694
rect 1996 3554 2036 3594
rect 1996 3454 2036 3494
rect 2140 3754 2180 3794
rect 2140 3654 2180 3694
rect 2140 3554 2180 3594
rect 2140 3454 2180 3494
rect 2428 3754 2468 3794
rect 2428 3654 2468 3694
rect 2428 3554 2468 3594
rect 2428 3454 2468 3494
rect 2572 3754 2612 3794
rect 2572 3654 2612 3694
rect 2572 3554 2612 3594
rect 2572 3454 2612 3494
rect 2716 3754 2756 3794
rect 2716 3654 2756 3694
rect 2716 3554 2756 3594
rect 2716 3454 2756 3494
rect 3004 3754 3044 3794
rect 3004 3654 3044 3694
rect 3004 3554 3044 3594
rect 3004 3454 3044 3494
rect 3148 3754 3188 3794
rect 3148 3654 3188 3694
rect 3148 3554 3188 3594
rect 3148 3454 3188 3494
rect 3292 3754 3332 3794
rect 4156 3754 4196 3794
rect 3292 3654 3332 3694
rect 3292 3554 3332 3594
rect 4156 3654 4196 3694
rect 4156 3554 4196 3594
rect 3292 3454 3332 3494
rect 4156 3454 4196 3494
rect 4300 3754 4340 3794
rect 4300 3654 4340 3694
rect 4300 3554 4340 3594
rect 4300 3454 4340 3494
rect 4444 3754 4484 3794
rect 4444 3654 4484 3694
rect 4444 3554 4484 3594
rect 4444 3454 4484 3494
rect 4732 3754 4772 3794
rect 4732 3654 4772 3694
rect 4732 3554 4772 3594
rect 4732 3454 4772 3494
rect 4876 3754 4916 3794
rect 4876 3654 4916 3694
rect 4876 3554 4916 3594
rect 4876 3454 4916 3494
rect 5020 3754 5060 3794
rect 5020 3654 5060 3694
rect 5020 3554 5060 3594
rect 5020 3454 5060 3494
rect 5308 3754 5348 3794
rect 5308 3654 5348 3694
rect 5308 3554 5348 3594
rect 5308 3454 5348 3494
rect 5452 3754 5492 3794
rect 5452 3654 5492 3694
rect 5452 3554 5492 3594
rect 5452 3454 5492 3494
rect 5596 3754 5636 3794
rect 5596 3654 5636 3694
rect 5596 3554 5636 3594
rect 5596 3454 5636 3494
rect 5884 3754 5924 3794
rect 5884 3654 5924 3694
rect 5884 3554 5924 3594
rect 5884 3454 5924 3494
rect 6028 3754 6068 3794
rect 6028 3654 6068 3694
rect 6028 3554 6068 3594
rect 6028 3454 6068 3494
rect 6172 3754 6212 3794
rect 6172 3654 6212 3694
rect 6172 3554 6212 3594
rect 6172 3454 6212 3494
rect 6460 3754 6500 3794
rect 6460 3654 6500 3694
rect 6460 3554 6500 3594
rect 6460 3454 6500 3494
rect 6604 3754 6644 3794
rect 6604 3654 6644 3694
rect 6604 3554 6644 3594
rect 6604 3454 6644 3494
rect 6748 3754 6788 3794
rect 7612 3754 7652 3794
rect 6748 3654 6788 3694
rect 6748 3554 6788 3594
rect 7612 3654 7652 3694
rect 7612 3554 7652 3594
rect 6748 3454 6788 3494
rect 7612 3454 7652 3494
rect 7756 3754 7796 3794
rect 7756 3654 7796 3694
rect 7756 3554 7796 3594
rect 7756 3454 7796 3494
rect 7900 3754 7940 3794
rect 7900 3654 7940 3694
rect 7900 3554 7940 3594
rect 7900 3454 7940 3494
rect 8188 3754 8228 3794
rect 8188 3654 8228 3694
rect 8188 3554 8228 3594
rect 8188 3454 8228 3494
rect 8332 3754 8372 3794
rect 8332 3654 8372 3694
rect 8332 3554 8372 3594
rect 8332 3454 8372 3494
rect 8476 3754 8516 3794
rect 8476 3654 8516 3694
rect 8476 3554 8516 3594
rect 8476 3454 8516 3494
rect 8764 3754 8804 3794
rect 8764 3654 8804 3694
rect 8764 3554 8804 3594
rect 8764 3454 8804 3494
rect 8908 3754 8948 3794
rect 8908 3654 8948 3694
rect 8908 3554 8948 3594
rect 8908 3454 8948 3494
rect 9052 3754 9092 3794
rect 9052 3654 9092 3694
rect 9052 3554 9092 3594
rect 9052 3454 9092 3494
rect 9340 3754 9380 3794
rect 9340 3654 9380 3694
rect 9340 3554 9380 3594
rect 9340 3454 9380 3494
rect 9484 3754 9524 3794
rect 9484 3654 9524 3694
rect 9484 3554 9524 3594
rect 9484 3454 9524 3494
rect 9628 3754 9668 3794
rect 9628 3654 9668 3694
rect 9628 3554 9668 3594
rect 9628 3454 9668 3494
rect 10204 3754 10244 3794
rect 10204 3654 10244 3694
rect 10204 3554 10244 3594
rect 10204 3454 10244 3494
rect 10348 3754 10388 3794
rect 10348 3654 10388 3694
rect 10348 3554 10388 3594
rect 10348 3454 10388 3494
rect 10492 3754 10532 3794
rect 10492 3654 10532 3694
rect 10492 3554 10532 3594
rect 10492 3454 10532 3494
rect 10780 3754 10820 3794
rect 10780 3654 10820 3694
rect 10780 3554 10820 3594
rect 10780 3454 10820 3494
rect 10924 3754 10964 3794
rect 10924 3654 10964 3694
rect 10924 3554 10964 3594
rect 10924 3454 10964 3494
rect 11068 3754 11108 3794
rect 11932 3754 11972 3794
rect 11068 3654 11108 3694
rect 11068 3554 11108 3594
rect 11932 3654 11972 3694
rect 11932 3554 11972 3594
rect 11068 3454 11108 3494
rect 11932 3454 11972 3494
rect 12076 3754 12116 3794
rect 12076 3654 12116 3694
rect 12076 3554 12116 3594
rect 12076 3454 12116 3494
rect 12220 3754 12260 3794
rect 12220 3654 12260 3694
rect 12220 3554 12260 3594
rect 12220 3454 12260 3494
rect 12508 3754 12548 3794
rect 12508 3654 12548 3694
rect 12508 3554 12548 3594
rect 12508 3454 12548 3494
rect 12652 3754 12692 3794
rect 12652 3654 12692 3694
rect 12652 3554 12692 3594
rect 12652 3454 12692 3494
rect 12796 3754 12836 3794
rect 12796 3654 12836 3694
rect 12796 3554 12836 3594
rect 12796 3454 12836 3494
rect 13660 3754 13700 3794
rect 13660 3654 13700 3694
rect 13660 3554 13700 3594
rect 13660 3454 13700 3494
rect 13804 3754 13844 3794
rect 13804 3654 13844 3694
rect 13804 3554 13844 3594
rect 13804 3454 13844 3494
rect 13948 3754 13988 3794
rect 13948 3654 13988 3694
rect 13948 3554 13988 3594
rect 13948 3454 13988 3494
rect 14236 3754 14276 3794
rect 14236 3654 14276 3694
rect 14236 3554 14276 3594
rect 14236 3454 14276 3494
rect 14380 3754 14420 3794
rect 14380 3654 14420 3694
rect 14380 3554 14420 3594
rect 14380 3454 14420 3494
rect 14524 3754 14564 3794
rect 14524 3654 14564 3694
rect 14524 3554 14564 3594
rect 14524 3454 14564 3494
rect 14812 3754 14852 3794
rect 14812 3654 14852 3694
rect 14812 3554 14852 3594
rect 14812 3454 14852 3494
rect 14956 3754 14996 3794
rect 14956 3654 14996 3694
rect 14956 3554 14996 3594
rect 14956 3454 14996 3494
rect 15100 3754 15140 3794
rect 16540 3754 16580 3794
rect 15100 3654 15140 3694
rect 15100 3554 15140 3594
rect 16540 3654 16580 3694
rect 16540 3554 16580 3594
rect 15100 3454 15140 3494
rect 16540 3454 16580 3494
rect 16684 3754 16724 3794
rect 16684 3654 16724 3694
rect 16684 3554 16724 3594
rect 16684 3454 16724 3494
rect 16828 3754 16868 3794
rect 16828 3654 16868 3694
rect 16828 3554 16868 3594
rect 16828 3454 16868 3494
rect 16972 3754 17012 3794
rect 16972 3654 17012 3694
rect 16972 3554 17012 3594
rect 16972 3454 17012 3494
rect 17116 3754 17156 3794
rect 17116 3654 17156 3694
rect 17116 3554 17156 3594
rect 17116 3454 17156 3494
rect 17260 3754 17300 3794
rect 17260 3654 17300 3694
rect 17260 3554 17300 3594
rect 17260 3454 17300 3494
rect 17404 3754 17444 3794
rect 17404 3654 17444 3694
rect 17404 3554 17444 3594
rect 17404 3454 17444 3494
rect 17548 3754 17588 3794
rect 17548 3654 17588 3694
rect 17548 3554 17588 3594
rect 17548 3454 17588 3494
rect 17692 3754 17732 3794
rect 17692 3654 17732 3694
rect 17692 3554 17732 3594
rect 17692 3454 17732 3494
rect 17836 3754 17876 3794
rect 17836 3654 17876 3694
rect 17836 3554 17876 3594
rect 17836 3454 17876 3494
rect 17980 3754 18020 3794
rect 17980 3654 18020 3694
rect 17980 3554 18020 3594
rect 17980 3454 18020 3494
rect 18124 3754 18164 3794
rect 18124 3654 18164 3694
rect 18124 3554 18164 3594
rect 18124 3454 18164 3494
rect 18268 3754 18308 3794
rect 18268 3654 18308 3694
rect 18268 3554 18308 3594
rect 18268 3454 18308 3494
rect 18412 3754 18452 3794
rect 18412 3654 18452 3694
rect 18412 3554 18452 3594
rect 18412 3454 18452 3494
rect 18556 3754 18596 3794
rect 18556 3654 18596 3694
rect 18556 3554 18596 3594
rect 18556 3454 18596 3494
rect 18700 3754 18740 3794
rect 18700 3654 18740 3694
rect 18700 3554 18740 3594
rect 18700 3454 18740 3494
rect 18844 3754 18884 3794
rect 18844 3654 18884 3694
rect 18844 3554 18884 3594
rect 18844 3454 18884 3494
rect 18988 3754 19028 3794
rect 18988 3654 19028 3694
rect 18988 3554 19028 3594
rect 18988 3454 19028 3494
rect 19132 3754 19172 3794
rect 19132 3654 19172 3694
rect 19132 3554 19172 3594
rect 19132 3454 19172 3494
rect 19276 3754 19316 3794
rect 19276 3654 19316 3694
rect 19276 3554 19316 3594
rect 19276 3454 19316 3494
rect 19420 3754 19460 3794
rect 19420 3654 19460 3694
rect 19420 3554 19460 3594
rect 19420 3454 19460 3494
rect 19564 3754 19604 3794
rect 19564 3654 19604 3694
rect 19564 3554 19604 3594
rect 19564 3454 19604 3494
rect 19708 3754 19748 3794
rect 19708 3654 19748 3694
rect 19708 3554 19748 3594
rect 19708 3454 19748 3494
rect 19852 3754 19892 3794
rect 19852 3654 19892 3694
rect 19852 3554 19892 3594
rect 19852 3454 19892 3494
rect 19996 3754 20036 3794
rect 19996 3654 20036 3694
rect 19996 3554 20036 3594
rect 19996 3454 20036 3494
rect 700 538 740 578
rect 700 438 740 478
rect 700 338 740 378
rect 700 238 740 278
rect 844 538 884 578
rect 844 438 884 478
rect 844 338 884 378
rect 844 238 884 278
rect 988 538 1028 578
rect 988 438 1028 478
rect 988 338 1028 378
rect 988 238 1028 278
rect 1276 538 1316 578
rect 1276 438 1316 478
rect 1276 338 1316 378
rect 1276 238 1316 278
rect 1420 538 1460 578
rect 1420 438 1460 478
rect 1420 338 1460 378
rect 1420 238 1460 278
rect 1564 538 1604 578
rect 1564 438 1604 478
rect 1564 338 1604 378
rect 1564 238 1604 278
rect 1852 538 1892 578
rect 1852 438 1892 478
rect 1852 338 1892 378
rect 1852 238 1892 278
rect 1996 538 2036 578
rect 1996 438 2036 478
rect 1996 338 2036 378
rect 1996 238 2036 278
rect 2140 538 2180 578
rect 2140 438 2180 478
rect 2140 338 2180 378
rect 2140 238 2180 278
rect 3004 538 3044 578
rect 3004 438 3044 478
rect 3004 338 3044 378
rect 3004 238 3044 278
rect 3148 538 3188 578
rect 3148 438 3188 478
rect 3148 338 3188 378
rect 3148 238 3188 278
rect 3292 538 3332 578
rect 3292 438 3332 478
rect 3292 338 3332 378
rect 3292 238 3332 278
rect 3580 538 3620 578
rect 3580 438 3620 478
rect 3580 338 3620 378
rect 3580 238 3620 278
rect 3724 538 3764 578
rect 3724 438 3764 478
rect 3724 338 3764 378
rect 3724 238 3764 278
rect 3868 538 3908 578
rect 3868 438 3908 478
rect 3868 338 3908 378
rect 3868 238 3908 278
rect 4156 538 4196 578
rect 4156 438 4196 478
rect 4156 338 4196 378
rect 4156 238 4196 278
rect 4300 538 4340 578
rect 4300 438 4340 478
rect 4300 338 4340 378
rect 4300 238 4340 278
rect 4444 538 4484 578
rect 5884 538 5924 578
rect 4444 438 4484 478
rect 4444 338 4484 378
rect 5884 438 5924 478
rect 5884 338 5924 378
rect 4444 238 4484 278
rect 5884 238 5924 278
rect 6028 538 6068 578
rect 6028 438 6068 478
rect 6028 338 6068 378
rect 6028 238 6068 278
rect 6172 538 6212 578
rect 6172 438 6212 478
rect 6172 338 6212 378
rect 6172 238 6212 278
rect 6460 538 6500 578
rect 6460 438 6500 478
rect 6460 338 6500 378
rect 6460 238 6500 278
rect 6604 538 6644 578
rect 6604 438 6644 478
rect 6604 338 6644 378
rect 6604 238 6644 278
rect 6748 538 6788 578
rect 6748 438 6788 478
rect 6748 338 6788 378
rect 6748 238 6788 278
rect 7036 538 7076 578
rect 7036 438 7076 478
rect 7036 338 7076 378
rect 7036 238 7076 278
rect 7180 538 7220 578
rect 7180 438 7220 478
rect 7180 338 7220 378
rect 7180 238 7220 278
rect 7324 538 7364 578
rect 7324 438 7364 478
rect 7324 338 7364 378
rect 7324 238 7364 278
rect 7612 538 7652 578
rect 7612 438 7652 478
rect 7612 338 7652 378
rect 7612 238 7652 278
rect 7756 538 7796 578
rect 7756 438 7796 478
rect 7756 338 7796 378
rect 7756 238 7796 278
rect 7900 538 7940 578
rect 7900 438 7940 478
rect 7900 338 7940 378
rect 7900 238 7940 278
rect 8188 538 8228 578
rect 8188 438 8228 478
rect 8188 338 8228 378
rect 8188 238 8228 278
rect 8332 538 8372 578
rect 8332 438 8372 478
rect 8332 338 8372 378
rect 8332 238 8372 278
rect 8476 538 8516 578
rect 9340 538 9380 578
rect 8476 438 8516 478
rect 8476 338 8516 378
rect 9340 438 9380 478
rect 9340 338 9380 378
rect 8476 238 8516 278
rect 9340 238 9380 278
rect 9484 538 9524 578
rect 9484 438 9524 478
rect 9484 338 9524 378
rect 9484 238 9524 278
rect 9628 538 9668 578
rect 9628 438 9668 478
rect 9628 338 9668 378
rect 9628 238 9668 278
rect 9916 538 9956 578
rect 9916 438 9956 478
rect 9916 338 9956 378
rect 9916 238 9956 278
rect 10060 538 10100 578
rect 10060 438 10100 478
rect 10060 338 10100 378
rect 10060 238 10100 278
rect 10204 538 10244 578
rect 10204 438 10244 478
rect 10204 338 10244 378
rect 10204 238 10244 278
rect 10492 538 10532 578
rect 10492 438 10532 478
rect 10492 338 10532 378
rect 10492 238 10532 278
rect 10636 538 10676 578
rect 10636 438 10676 478
rect 10636 338 10676 378
rect 10636 238 10676 278
rect 10780 538 10820 578
rect 10780 438 10820 478
rect 10780 338 10820 378
rect 10780 238 10820 278
rect 11068 538 11108 578
rect 11068 438 11108 478
rect 11068 338 11108 378
rect 11068 238 11108 278
rect 11212 538 11252 578
rect 11212 438 11252 478
rect 11212 338 11252 378
rect 11212 238 11252 278
rect 11356 538 11396 578
rect 11356 438 11396 478
rect 11356 338 11396 378
rect 11356 238 11396 278
rect 11932 538 11972 578
rect 11932 438 11972 478
rect 11932 338 11972 378
rect 11932 238 11972 278
rect 12076 538 12116 578
rect 12076 438 12116 478
rect 12076 338 12116 378
rect 12076 238 12116 278
rect 12220 538 12260 578
rect 12220 438 12260 478
rect 12220 338 12260 378
rect 12220 238 12260 278
rect 12508 538 12548 578
rect 12508 438 12548 478
rect 12508 338 12548 378
rect 12508 238 12548 278
rect 12652 538 12692 578
rect 12652 438 12692 478
rect 12652 338 12692 378
rect 12652 238 12692 278
rect 12796 538 12836 578
rect 12796 438 12836 478
rect 12796 338 12836 378
rect 12796 238 12836 278
rect 13084 538 13124 578
rect 13084 438 13124 478
rect 13084 338 13124 378
rect 13084 238 13124 278
rect 13228 538 13268 578
rect 13228 438 13268 478
rect 13228 338 13268 378
rect 13228 238 13268 278
rect 13372 538 13412 578
rect 13372 438 13412 478
rect 13372 338 13412 378
rect 13372 238 13412 278
rect 13660 538 13700 578
rect 13660 438 13700 478
rect 13660 338 13700 378
rect 13660 238 13700 278
rect 13804 538 13844 578
rect 13804 438 13844 478
rect 13804 338 13844 378
rect 13804 238 13844 278
rect 13948 538 13988 578
rect 14812 538 14852 578
rect 13948 438 13988 478
rect 13948 338 13988 378
rect 14812 438 14852 478
rect 14812 338 14852 378
rect 13948 238 13988 278
rect 14812 238 14852 278
rect 14956 538 14996 578
rect 14956 438 14996 478
rect 14956 338 14996 378
rect 14956 238 14996 278
rect 15100 538 15140 578
rect 15100 438 15140 478
rect 15100 338 15140 378
rect 15100 238 15140 278
rect 15388 538 15428 578
rect 15388 438 15428 478
rect 15388 338 15428 378
rect 15388 238 15428 278
rect 15532 538 15572 578
rect 15532 438 15572 478
rect 15532 338 15572 378
rect 15532 238 15572 278
rect 15676 538 15716 578
rect 15676 438 15716 478
rect 15676 338 15716 378
rect 15676 238 15716 278
rect 15964 538 16004 578
rect 15964 438 16004 478
rect 15964 338 16004 378
rect 15964 238 16004 278
rect 16108 538 16148 578
rect 16108 438 16148 478
rect 16108 338 16148 378
rect 16108 238 16148 278
rect 16252 538 16292 578
rect 16252 438 16292 478
rect 16252 338 16292 378
rect 16252 238 16292 278
rect 16396 538 16436 578
rect 16396 438 16436 478
rect 16396 338 16436 378
rect 16396 238 16436 278
rect 16540 538 16580 578
rect 17404 538 17444 578
rect 16540 438 16580 478
rect 16540 338 16580 378
rect 17404 438 17444 478
rect 17404 338 17444 378
rect 16540 238 16580 278
rect 17404 238 17444 278
rect 17548 538 17588 578
rect 17548 438 17588 478
rect 17548 338 17588 378
rect 17548 238 17588 278
rect 17692 538 17732 578
rect 17692 438 17732 478
rect 17692 338 17732 378
rect 17692 238 17732 278
rect 17836 538 17876 578
rect 17836 438 17876 478
rect 17836 338 17876 378
rect 17836 238 17876 278
rect 17980 538 18020 578
rect 17980 438 18020 478
rect 17980 338 18020 378
rect 17980 238 18020 278
rect 18124 538 18164 578
rect 18124 438 18164 478
rect 18124 338 18164 378
rect 18124 238 18164 278
rect 18268 538 18308 578
rect 18268 438 18308 478
rect 18268 338 18308 378
rect 18268 238 18308 278
rect 18412 538 18452 578
rect 18412 438 18452 478
rect 18412 338 18452 378
rect 18412 238 18452 278
rect 18556 538 18596 578
rect 18556 438 18596 478
rect 18556 338 18596 378
rect 18556 238 18596 278
rect 18700 538 18740 578
rect 18700 438 18740 478
rect 18700 338 18740 378
rect 18700 238 18740 278
rect 18844 538 18884 578
rect 18844 438 18884 478
rect 18844 338 18884 378
rect 18844 238 18884 278
rect 18988 538 19028 578
rect 18988 438 19028 478
rect 18988 338 19028 378
rect 18988 238 19028 278
rect 19132 538 19172 578
rect 19132 438 19172 478
rect 19132 338 19172 378
rect 19132 238 19172 278
rect 19276 538 19316 578
rect 19276 438 19316 478
rect 19276 338 19316 378
rect 19276 238 19316 278
rect 19420 538 19460 578
rect 19420 438 19460 478
rect 19420 338 19460 378
rect 19420 238 19460 278
rect 19564 538 19604 578
rect 19564 438 19604 478
rect 19564 338 19604 378
rect 19564 238 19604 278
rect 19708 538 19748 578
rect 19708 438 19748 478
rect 19708 338 19748 378
rect 19708 238 19748 278
rect 19852 538 19892 578
rect 19852 438 19892 478
rect 19852 338 19892 378
rect 19852 238 19892 278
rect 19996 538 20036 578
rect 19996 438 20036 478
rect 19996 338 20036 378
rect 19996 238 20036 278
rect 20140 538 20180 578
rect 20140 438 20180 478
rect 20140 338 20180 378
rect 20140 238 20180 278
rect 20284 538 20324 578
rect 20284 438 20324 478
rect 20284 338 20324 378
rect 20284 238 20324 278
rect 20428 538 20468 578
rect 20428 438 20468 478
rect 20428 338 20468 378
rect 20428 238 20468 278
rect 20572 538 20612 578
rect 20572 438 20612 478
rect 20572 338 20612 378
rect 20572 238 20612 278
rect 20716 538 20756 578
rect 20716 438 20756 478
rect 20716 338 20756 378
rect 20716 238 20756 278
rect 20860 538 20900 578
rect 20860 438 20900 478
rect 20860 338 20900 378
rect 20860 238 20900 278
<< psubdiff >>
rect 114 2588 462 2630
rect 114 2500 124 2588
rect 164 2500 268 2588
rect 308 2500 412 2588
rect 452 2500 462 2588
rect 114 2458 462 2500
rect 3570 2588 3918 2630
rect 3570 2500 3580 2588
rect 3620 2500 3724 2588
rect 3764 2500 3868 2588
rect 3908 2500 3918 2588
rect 3570 2458 3918 2500
rect 7026 2588 7374 2630
rect 7026 2500 7036 2588
rect 7076 2500 7180 2588
rect 7220 2500 7324 2588
rect 7364 2500 7374 2588
rect 7026 2458 7374 2500
rect 11346 2588 11694 2630
rect 11346 2500 11356 2588
rect 11396 2500 11500 2588
rect 11540 2500 11644 2588
rect 11684 2500 11694 2588
rect 11346 2458 11694 2500
rect 15378 2588 15726 2630
rect 15378 2500 15388 2588
rect 15428 2500 15532 2588
rect 15572 2500 15676 2588
rect 15716 2500 15726 2588
rect 15378 2458 15726 2500
rect 15954 2588 16302 2630
rect 15954 2500 15964 2588
rect 16004 2500 16108 2588
rect 16148 2500 16252 2588
rect 16292 2500 16302 2588
rect 15954 2458 16302 2500
rect 114 1532 462 1574
rect 114 1444 124 1532
rect 164 1444 268 1532
rect 308 1444 412 1532
rect 452 1444 462 1532
rect 114 1402 462 1444
rect 4722 1532 5070 1574
rect 4722 1444 4732 1532
rect 4772 1444 4876 1532
rect 4916 1444 5020 1532
rect 5060 1444 5070 1532
rect 4722 1402 5070 1444
rect 5298 1532 5646 1574
rect 5298 1444 5308 1532
rect 5348 1444 5452 1532
rect 5492 1444 5596 1532
rect 5636 1444 5646 1532
rect 5298 1402 5646 1444
rect 8754 1532 9102 1574
rect 8754 1444 8764 1532
rect 8804 1444 8908 1532
rect 8948 1444 9052 1532
rect 9092 1444 9102 1532
rect 8754 1402 9102 1444
rect 14226 1532 14574 1574
rect 14226 1444 14236 1532
rect 14276 1444 14380 1532
rect 14420 1444 14524 1532
rect 14564 1444 14574 1532
rect 14226 1402 14574 1444
rect 16818 1532 17166 1574
rect 16818 1444 16828 1532
rect 16868 1444 16972 1532
rect 17012 1444 17116 1532
rect 17156 1444 17166 1532
rect 16818 1402 17166 1444
<< nsubdiff >>
rect 114 3704 462 3728
rect 114 3552 124 3704
rect 164 3552 268 3704
rect 308 3552 412 3704
rect 452 3552 462 3704
rect 114 3528 462 3552
rect 3570 3704 3918 3728
rect 3570 3552 3580 3704
rect 3620 3552 3724 3704
rect 3764 3552 3868 3704
rect 3908 3552 3918 3704
rect 3570 3528 3918 3552
rect 7026 3704 7374 3728
rect 7026 3552 7036 3704
rect 7076 3552 7180 3704
rect 7220 3552 7324 3704
rect 7364 3552 7374 3704
rect 7026 3528 7374 3552
rect 11346 3704 11694 3728
rect 11346 3552 11356 3704
rect 11396 3552 11500 3704
rect 11540 3552 11644 3704
rect 11684 3552 11694 3704
rect 11346 3528 11694 3552
rect 15378 3704 15726 3728
rect 15378 3552 15388 3704
rect 15428 3552 15532 3704
rect 15572 3552 15676 3704
rect 15716 3552 15726 3704
rect 15378 3528 15726 3552
rect 15954 3704 16302 3728
rect 15954 3552 15964 3704
rect 16004 3552 16108 3704
rect 16148 3552 16252 3704
rect 16292 3552 16302 3704
rect 15954 3528 16302 3552
rect 114 480 462 504
rect 114 328 124 480
rect 164 328 268 480
rect 308 328 412 480
rect 452 328 462 480
rect 114 304 462 328
rect 4722 480 5070 504
rect 4722 328 4732 480
rect 4772 328 4876 480
rect 4916 328 5020 480
rect 5060 328 5070 480
rect 4722 304 5070 328
rect 5298 480 5646 504
rect 5298 328 5308 480
rect 5348 328 5452 480
rect 5492 328 5596 480
rect 5636 328 5646 480
rect 5298 304 5646 328
rect 8754 480 9102 504
rect 8754 328 8764 480
rect 8804 328 8908 480
rect 8948 328 9052 480
rect 9092 328 9102 480
rect 8754 304 9102 328
rect 14226 480 14574 504
rect 14226 328 14236 480
rect 14276 328 14380 480
rect 14420 328 14524 480
rect 14564 328 14574 480
rect 14226 304 14574 328
rect 16818 480 17166 504
rect 16818 328 16828 480
rect 16868 328 16972 480
rect 17012 328 17116 480
rect 17156 328 17166 480
rect 16818 304 17166 328
<< psubdiffcont >>
rect 124 2500 164 2588
rect 268 2500 308 2588
rect 412 2500 452 2588
rect 3580 2500 3620 2588
rect 3724 2500 3764 2588
rect 3868 2500 3908 2588
rect 7036 2500 7076 2588
rect 7180 2500 7220 2588
rect 7324 2500 7364 2588
rect 11356 2500 11396 2588
rect 11500 2500 11540 2588
rect 11644 2500 11684 2588
rect 15388 2500 15428 2588
rect 15532 2500 15572 2588
rect 15676 2500 15716 2588
rect 15964 2500 16004 2588
rect 16108 2500 16148 2588
rect 16252 2500 16292 2588
rect 124 1444 164 1532
rect 268 1444 308 1532
rect 412 1444 452 1532
rect 4732 1444 4772 1532
rect 4876 1444 4916 1532
rect 5020 1444 5060 1532
rect 5308 1444 5348 1532
rect 5452 1444 5492 1532
rect 5596 1444 5636 1532
rect 8764 1444 8804 1532
rect 8908 1444 8948 1532
rect 9052 1444 9092 1532
rect 14236 1444 14276 1532
rect 14380 1444 14420 1532
rect 14524 1444 14564 1532
rect 16828 1444 16868 1532
rect 16972 1444 17012 1532
rect 17116 1444 17156 1532
<< nsubdiffcont >>
rect 124 3552 164 3704
rect 268 3552 308 3704
rect 412 3552 452 3704
rect 3580 3552 3620 3704
rect 3724 3552 3764 3704
rect 3868 3552 3908 3704
rect 7036 3552 7076 3704
rect 7180 3552 7220 3704
rect 7324 3552 7364 3704
rect 11356 3552 11396 3704
rect 11500 3552 11540 3704
rect 11644 3552 11684 3704
rect 15388 3552 15428 3704
rect 15532 3552 15572 3704
rect 15676 3552 15716 3704
rect 15964 3552 16004 3704
rect 16108 3552 16148 3704
rect 16252 3552 16292 3704
rect 124 328 164 480
rect 268 328 308 480
rect 412 328 452 480
rect 4732 328 4772 480
rect 4876 328 4916 480
rect 5020 328 5060 480
rect 5308 328 5348 480
rect 5452 328 5492 480
rect 5596 328 5636 480
rect 8764 328 8804 480
rect 8908 328 8948 480
rect 9052 328 9092 480
rect 14236 328 14276 480
rect 14380 328 14420 480
rect 14524 328 14564 480
rect 16828 328 16868 480
rect 16972 328 17012 480
rect 17116 328 17156 480
<< poly >>
rect 778 3864 808 3900
rect 922 3864 952 3900
rect 1354 3864 1384 3900
rect 1498 3864 1528 3900
rect 1930 3864 1960 3900
rect 2074 3864 2104 3900
rect 2506 3864 2536 3900
rect 2650 3864 2680 3900
rect 3080 3864 3110 3900
rect 3224 3864 3254 3900
rect 4232 3864 4262 3900
rect 4376 3864 4406 3900
rect 4808 3864 4838 3900
rect 4952 3864 4982 3900
rect 5384 3864 5414 3900
rect 5528 3864 5558 3900
rect 5960 3864 5990 3900
rect 6104 3864 6134 3900
rect 6536 3864 6566 3900
rect 6680 3864 6710 3900
rect 7688 3864 7718 3900
rect 7832 3864 7862 3900
rect 8264 3864 8294 3900
rect 8408 3864 8438 3900
rect 8840 3864 8870 3900
rect 8984 3864 9014 3900
rect 9416 3864 9446 3900
rect 9560 3864 9590 3900
rect 10280 3864 10310 3900
rect 10424 3864 10454 3900
rect 10856 3864 10886 3900
rect 11000 3864 11030 3900
rect 12008 3864 12038 3900
rect 12152 3864 12182 3900
rect 12584 3864 12614 3900
rect 12728 3864 12758 3900
rect 13736 3864 13766 3900
rect 13880 3864 13910 3900
rect 14312 3864 14342 3900
rect 14456 3864 14486 3900
rect 14888 3864 14918 3900
rect 15032 3864 15062 3900
rect 16618 3864 16648 3900
rect 16762 3864 16792 3900
rect 16906 3864 16936 3900
rect 17050 3864 17080 3900
rect 17194 3864 17224 3900
rect 17338 3864 17368 3900
rect 17482 3864 17512 3900
rect 17626 3864 17656 3900
rect 17770 3864 17800 3900
rect 17914 3864 17944 3900
rect 18058 3864 18088 3900
rect 18202 3864 18232 3900
rect 18346 3864 18376 3900
rect 18490 3864 18520 3900
rect 18634 3864 18664 3900
rect 18778 3864 18808 3900
rect 18922 3864 18952 3900
rect 19066 3864 19096 3900
rect 19210 3864 19240 3900
rect 19354 3864 19384 3900
rect 19498 3864 19528 3900
rect 19642 3864 19672 3900
rect 19786 3864 19816 3900
rect 19930 3864 19960 3900
rect 778 3348 808 3384
rect 922 3348 952 3384
rect 778 3329 952 3348
rect 778 3295 790 3329
rect 824 3295 898 3329
rect 932 3295 952 3329
rect 778 3276 952 3295
rect 1354 3348 1384 3384
rect 1498 3348 1528 3384
rect 1354 3329 1528 3348
rect 1354 3295 1366 3329
rect 1400 3295 1474 3329
rect 1508 3295 1528 3329
rect 1354 3276 1528 3295
rect 1930 3348 1960 3384
rect 2074 3348 2104 3384
rect 1930 3329 2104 3348
rect 1930 3295 1942 3329
rect 1976 3295 2050 3329
rect 2084 3295 2104 3329
rect 1930 3276 2104 3295
rect 2506 3348 2536 3384
rect 2650 3348 2680 3384
rect 2506 3329 2680 3348
rect 2506 3295 2518 3329
rect 2552 3295 2626 3329
rect 2660 3295 2680 3329
rect 2506 3276 2680 3295
rect 3080 3348 3110 3384
rect 3224 3348 3254 3384
rect 3080 3329 3254 3348
rect 3080 3295 3100 3329
rect 3134 3295 3208 3329
rect 3242 3295 3254 3329
rect 3080 3276 3254 3295
rect 4232 3348 4262 3384
rect 4376 3348 4406 3384
rect 4232 3329 4406 3348
rect 4232 3295 4252 3329
rect 4286 3295 4360 3329
rect 4394 3295 4406 3329
rect 4232 3276 4406 3295
rect 4808 3348 4838 3384
rect 4952 3348 4982 3384
rect 4808 3329 4982 3348
rect 4808 3295 4828 3329
rect 4862 3295 4936 3329
rect 4970 3295 4982 3329
rect 4808 3276 4982 3295
rect 5384 3348 5414 3384
rect 5528 3348 5558 3384
rect 5384 3329 5558 3348
rect 5384 3295 5404 3329
rect 5438 3295 5512 3329
rect 5546 3295 5558 3329
rect 5384 3276 5558 3295
rect 5960 3348 5990 3384
rect 6104 3348 6134 3384
rect 6536 3348 6566 3384
rect 5960 3329 6134 3348
rect 5960 3295 5980 3329
rect 6014 3295 6088 3329
rect 6122 3295 6134 3329
rect 5960 3276 6134 3295
rect 6446 3330 6566 3348
rect 6446 3294 6468 3330
rect 6504 3294 6566 3330
rect 6446 3276 6566 3294
rect 6680 3348 6710 3384
rect 7688 3348 7718 3384
rect 7832 3348 7862 3384
rect 6680 3330 6800 3348
rect 6680 3294 6752 3330
rect 6788 3294 6800 3330
rect 6680 3276 6800 3294
rect 7688 3329 7862 3348
rect 7688 3295 7708 3329
rect 7742 3295 7816 3329
rect 7850 3295 7862 3329
rect 7688 3276 7862 3295
rect 8264 3348 8294 3384
rect 8408 3348 8438 3384
rect 8264 3329 8438 3348
rect 8264 3295 8284 3329
rect 8318 3295 8392 3329
rect 8426 3295 8438 3329
rect 8264 3276 8438 3295
rect 8840 3348 8870 3384
rect 8984 3348 9014 3384
rect 9416 3348 9446 3384
rect 8840 3329 9014 3348
rect 8840 3295 8860 3329
rect 8894 3295 8968 3329
rect 9002 3295 9014 3329
rect 8840 3276 9014 3295
rect 9326 3330 9446 3348
rect 9326 3294 9348 3330
rect 9384 3294 9446 3330
rect 9326 3276 9446 3294
rect 9560 3348 9590 3384
rect 10280 3348 10310 3384
rect 10424 3348 10454 3384
rect 9560 3330 9680 3348
rect 9560 3294 9632 3330
rect 9668 3294 9680 3330
rect 9560 3276 9680 3294
rect 10280 3329 10454 3348
rect 10280 3295 10300 3329
rect 10334 3295 10408 3329
rect 10442 3295 10454 3329
rect 10280 3276 10454 3295
rect 10856 3348 10886 3384
rect 11000 3348 11030 3384
rect 10856 3329 11030 3348
rect 10856 3295 10876 3329
rect 10910 3295 10984 3329
rect 11018 3295 11030 3329
rect 10856 3276 11030 3295
rect 12008 3348 12038 3384
rect 12152 3348 12182 3384
rect 12008 3329 12182 3348
rect 12008 3295 12028 3329
rect 12062 3295 12136 3329
rect 12170 3295 12182 3329
rect 12008 3276 12182 3295
rect 12584 3348 12614 3384
rect 12728 3348 12758 3384
rect 12584 3329 12758 3348
rect 12584 3295 12604 3329
rect 12638 3295 12712 3329
rect 12746 3295 12758 3329
rect 12584 3276 12758 3295
rect 13736 3348 13766 3384
rect 13880 3348 13910 3384
rect 13736 3329 13910 3348
rect 13736 3295 13756 3329
rect 13790 3295 13864 3329
rect 13898 3295 13910 3329
rect 13736 3276 13910 3295
rect 14312 3348 14342 3384
rect 14456 3348 14486 3384
rect 14312 3329 14486 3348
rect 14312 3295 14332 3329
rect 14366 3295 14440 3329
rect 14474 3295 14486 3329
rect 14312 3276 14486 3295
rect 14888 3348 14918 3384
rect 15032 3348 15062 3384
rect 14888 3329 15062 3348
rect 14888 3295 14908 3329
rect 14942 3295 15016 3329
rect 15050 3295 15062 3329
rect 14888 3276 15062 3295
rect 16618 3348 16648 3384
rect 16762 3348 16792 3384
rect 16618 3329 16792 3348
rect 16618 3295 16630 3329
rect 16664 3295 16738 3329
rect 16772 3295 16792 3329
rect 16618 3276 16792 3295
rect 16906 3348 16936 3384
rect 17050 3348 17080 3384
rect 16906 3329 17080 3348
rect 16906 3295 16918 3329
rect 16952 3295 17026 3329
rect 17060 3295 17080 3329
rect 16906 3276 17080 3295
rect 17194 3348 17224 3384
rect 17338 3348 17368 3384
rect 17194 3329 17368 3348
rect 17194 3295 17206 3329
rect 17240 3295 17314 3329
rect 17348 3295 17368 3329
rect 17194 3276 17368 3295
rect 17482 3348 17512 3384
rect 17626 3348 17656 3384
rect 17482 3329 17656 3348
rect 17482 3295 17494 3329
rect 17528 3295 17602 3329
rect 17636 3295 17656 3329
rect 17482 3276 17656 3295
rect 17770 3348 17800 3384
rect 17914 3348 17944 3384
rect 17770 3329 17944 3348
rect 17770 3295 17782 3329
rect 17816 3295 17890 3329
rect 17924 3295 17944 3329
rect 17770 3276 17944 3295
rect 18058 3348 18088 3384
rect 18202 3348 18232 3384
rect 18058 3329 18232 3348
rect 18058 3295 18070 3329
rect 18104 3295 18178 3329
rect 18212 3295 18232 3329
rect 18058 3276 18232 3295
rect 18346 3348 18376 3384
rect 18490 3348 18520 3384
rect 18346 3329 18520 3348
rect 18346 3295 18358 3329
rect 18392 3295 18466 3329
rect 18500 3295 18520 3329
rect 18346 3276 18520 3295
rect 18634 3348 18664 3384
rect 18778 3348 18808 3384
rect 18634 3329 18808 3348
rect 18634 3295 18646 3329
rect 18680 3295 18754 3329
rect 18788 3295 18808 3329
rect 18634 3276 18808 3295
rect 18922 3348 18952 3384
rect 19066 3348 19096 3384
rect 18922 3329 19096 3348
rect 18922 3295 18934 3329
rect 18968 3295 19042 3329
rect 19076 3295 19096 3329
rect 18922 3276 19096 3295
rect 19210 3348 19240 3384
rect 19354 3348 19384 3384
rect 19210 3329 19384 3348
rect 19210 3295 19222 3329
rect 19256 3295 19330 3329
rect 19364 3295 19384 3329
rect 19210 3276 19384 3295
rect 19498 3348 19528 3384
rect 19642 3348 19672 3384
rect 19498 3329 19672 3348
rect 19498 3295 19510 3329
rect 19544 3295 19618 3329
rect 19652 3295 19672 3329
rect 19498 3276 19672 3295
rect 19786 3348 19816 3384
rect 19930 3348 19960 3384
rect 19786 3329 19960 3348
rect 19786 3295 19798 3329
rect 19832 3295 19906 3329
rect 19940 3295 19960 3329
rect 19786 3276 19960 3295
rect 778 2753 952 2772
rect 778 2719 790 2753
rect 824 2719 898 2753
rect 932 2719 952 2753
rect 778 2700 952 2719
rect 778 2664 808 2700
rect 922 2664 952 2700
rect 1354 2753 1528 2772
rect 1354 2719 1366 2753
rect 1400 2719 1474 2753
rect 1508 2719 1528 2753
rect 1354 2700 1528 2719
rect 1354 2664 1384 2700
rect 1498 2664 1528 2700
rect 1930 2753 2104 2772
rect 1930 2719 1942 2753
rect 1976 2719 2050 2753
rect 2084 2719 2104 2753
rect 1930 2700 2104 2719
rect 1930 2664 1960 2700
rect 2074 2664 2104 2700
rect 2506 2753 2680 2772
rect 2506 2719 2518 2753
rect 2552 2719 2626 2753
rect 2660 2719 2680 2753
rect 2506 2700 2680 2719
rect 2506 2664 2536 2700
rect 2650 2664 2680 2700
rect 3080 2753 3254 2772
rect 3080 2719 3100 2753
rect 3134 2719 3208 2753
rect 3242 2719 3254 2753
rect 3080 2700 3254 2719
rect 3080 2664 3110 2700
rect 3224 2664 3254 2700
rect 4232 2753 4406 2772
rect 4232 2719 4252 2753
rect 4286 2719 4360 2753
rect 4394 2719 4406 2753
rect 4232 2700 4406 2719
rect 4232 2664 4262 2700
rect 4376 2664 4406 2700
rect 4808 2753 4982 2772
rect 4808 2719 4828 2753
rect 4862 2719 4936 2753
rect 4970 2719 4982 2753
rect 4808 2700 4982 2719
rect 4808 2664 4838 2700
rect 4952 2664 4982 2700
rect 5384 2753 5558 2772
rect 5384 2719 5404 2753
rect 5438 2719 5512 2753
rect 5546 2719 5558 2753
rect 5384 2700 5558 2719
rect 5384 2664 5414 2700
rect 5528 2664 5558 2700
rect 5960 2753 6134 2772
rect 5960 2719 5980 2753
rect 6014 2719 6088 2753
rect 6122 2719 6134 2753
rect 5960 2700 6134 2719
rect 6446 2754 6566 2772
rect 6446 2718 6468 2754
rect 6504 2718 6566 2754
rect 6446 2700 6566 2718
rect 5960 2664 5990 2700
rect 6104 2664 6134 2700
rect 6536 2664 6566 2700
rect 6680 2754 6800 2772
rect 6680 2718 6746 2754
rect 6782 2718 6800 2754
rect 6680 2700 6800 2718
rect 7688 2753 7862 2772
rect 7688 2719 7708 2753
rect 7742 2719 7816 2753
rect 7850 2719 7862 2753
rect 7688 2700 7862 2719
rect 6680 2664 6710 2700
rect 7688 2664 7718 2700
rect 7832 2664 7862 2700
rect 8264 2753 8438 2772
rect 8264 2719 8284 2753
rect 8318 2719 8392 2753
rect 8426 2719 8438 2753
rect 8264 2700 8438 2719
rect 8264 2664 8294 2700
rect 8408 2664 8438 2700
rect 8840 2753 9014 2772
rect 8840 2719 8860 2753
rect 8894 2719 8968 2753
rect 9002 2719 9014 2753
rect 8840 2700 9014 2719
rect 9326 2754 9446 2772
rect 9326 2718 9348 2754
rect 9384 2718 9446 2754
rect 9326 2700 9446 2718
rect 8840 2664 8870 2700
rect 8984 2664 9014 2700
rect 9416 2664 9446 2700
rect 9560 2754 9680 2772
rect 9560 2718 9626 2754
rect 9662 2718 9680 2754
rect 9560 2700 9680 2718
rect 10280 2753 10454 2772
rect 10280 2719 10300 2753
rect 10334 2719 10408 2753
rect 10442 2719 10454 2753
rect 10280 2700 10454 2719
rect 9560 2664 9590 2700
rect 10280 2664 10310 2700
rect 10424 2664 10454 2700
rect 10856 2753 11030 2772
rect 10856 2719 10876 2753
rect 10910 2719 10984 2753
rect 11018 2719 11030 2753
rect 10856 2700 11030 2719
rect 10856 2664 10886 2700
rect 11000 2664 11030 2700
rect 12008 2753 12182 2772
rect 12008 2719 12028 2753
rect 12062 2719 12136 2753
rect 12170 2719 12182 2753
rect 12008 2700 12182 2719
rect 12008 2664 12038 2700
rect 12152 2664 12182 2700
rect 12584 2753 12758 2772
rect 12584 2719 12604 2753
rect 12638 2719 12712 2753
rect 12746 2719 12758 2753
rect 12584 2700 12758 2719
rect 12584 2664 12614 2700
rect 12728 2664 12758 2700
rect 13736 2753 13910 2772
rect 13736 2719 13756 2753
rect 13790 2719 13864 2753
rect 13898 2719 13910 2753
rect 13736 2700 13910 2719
rect 13736 2664 13766 2700
rect 13880 2664 13910 2700
rect 14312 2753 14486 2772
rect 14312 2719 14332 2753
rect 14366 2719 14440 2753
rect 14474 2719 14486 2753
rect 14312 2700 14486 2719
rect 14312 2664 14342 2700
rect 14456 2664 14486 2700
rect 14888 2753 15062 2772
rect 14888 2719 14908 2753
rect 14942 2719 15016 2753
rect 15050 2719 15062 2753
rect 14888 2700 15062 2719
rect 14888 2664 14918 2700
rect 15032 2664 15062 2700
rect 16618 2753 16792 2772
rect 16618 2719 16630 2753
rect 16664 2719 16738 2753
rect 16772 2719 16792 2753
rect 16618 2700 16792 2719
rect 16618 2664 16648 2700
rect 16762 2664 16792 2700
rect 16906 2753 17080 2772
rect 16906 2719 16918 2753
rect 16952 2719 17026 2753
rect 17060 2719 17080 2753
rect 16906 2700 17080 2719
rect 16906 2664 16936 2700
rect 17050 2664 17080 2700
rect 17194 2753 17368 2772
rect 17194 2719 17206 2753
rect 17240 2719 17314 2753
rect 17348 2719 17368 2753
rect 17194 2700 17368 2719
rect 17194 2664 17224 2700
rect 17338 2664 17368 2700
rect 17482 2753 17656 2772
rect 17482 2719 17494 2753
rect 17528 2719 17602 2753
rect 17636 2719 17656 2753
rect 17482 2700 17656 2719
rect 17482 2664 17512 2700
rect 17626 2664 17656 2700
rect 17770 2753 17944 2772
rect 17770 2719 17782 2753
rect 17816 2719 17890 2753
rect 17924 2719 17944 2753
rect 17770 2700 17944 2719
rect 17770 2664 17800 2700
rect 17914 2664 17944 2700
rect 18058 2753 18232 2772
rect 18058 2719 18070 2753
rect 18104 2719 18178 2753
rect 18212 2719 18232 2753
rect 18058 2700 18232 2719
rect 18058 2664 18088 2700
rect 18202 2664 18232 2700
rect 18346 2753 18520 2772
rect 18346 2719 18358 2753
rect 18392 2719 18466 2753
rect 18500 2719 18520 2753
rect 18346 2700 18520 2719
rect 18346 2664 18376 2700
rect 18490 2664 18520 2700
rect 18634 2753 18808 2772
rect 18634 2719 18646 2753
rect 18680 2719 18754 2753
rect 18788 2719 18808 2753
rect 18634 2700 18808 2719
rect 18634 2664 18664 2700
rect 18778 2664 18808 2700
rect 18922 2753 19096 2772
rect 18922 2719 18934 2753
rect 18968 2719 19042 2753
rect 19076 2719 19096 2753
rect 18922 2700 19096 2719
rect 18922 2664 18952 2700
rect 19066 2664 19096 2700
rect 19210 2753 19384 2772
rect 19210 2719 19222 2753
rect 19256 2719 19330 2753
rect 19364 2719 19384 2753
rect 19210 2700 19384 2719
rect 19210 2664 19240 2700
rect 19354 2664 19384 2700
rect 19498 2753 19672 2772
rect 19498 2719 19510 2753
rect 19544 2719 19618 2753
rect 19652 2719 19672 2753
rect 19498 2700 19672 2719
rect 19498 2664 19528 2700
rect 19642 2664 19672 2700
rect 19786 2753 19960 2772
rect 19786 2719 19798 2753
rect 19832 2719 19906 2753
rect 19940 2719 19960 2753
rect 19786 2700 19960 2719
rect 19786 2664 19816 2700
rect 19930 2664 19960 2700
rect 778 2388 808 2424
rect 922 2388 952 2424
rect 1354 2388 1384 2424
rect 1498 2388 1528 2424
rect 1930 2388 1960 2424
rect 2074 2388 2104 2424
rect 2506 2388 2536 2424
rect 2650 2388 2680 2424
rect 3080 2388 3110 2424
rect 3224 2388 3254 2424
rect 4232 2388 4262 2424
rect 4376 2388 4406 2424
rect 4808 2388 4838 2424
rect 4952 2388 4982 2424
rect 5384 2388 5414 2424
rect 5528 2388 5558 2424
rect 5960 2388 5990 2424
rect 6104 2388 6134 2424
rect 6536 2388 6566 2424
rect 6680 2388 6710 2424
rect 7688 2388 7718 2424
rect 7832 2388 7862 2424
rect 8264 2388 8294 2424
rect 8408 2388 8438 2424
rect 8840 2388 8870 2424
rect 8984 2388 9014 2424
rect 9416 2388 9446 2424
rect 9560 2388 9590 2424
rect 10280 2388 10310 2424
rect 10424 2388 10454 2424
rect 10856 2388 10886 2424
rect 11000 2388 11030 2424
rect 12008 2388 12038 2424
rect 12152 2388 12182 2424
rect 12584 2388 12614 2424
rect 12728 2388 12758 2424
rect 13736 2388 13766 2424
rect 13880 2388 13910 2424
rect 14312 2388 14342 2424
rect 14456 2388 14486 2424
rect 14888 2388 14918 2424
rect 15032 2388 15062 2424
rect 16618 2388 16648 2424
rect 16762 2388 16792 2424
rect 16906 2388 16936 2424
rect 17050 2388 17080 2424
rect 17194 2388 17224 2424
rect 17338 2388 17368 2424
rect 17482 2388 17512 2424
rect 17626 2388 17656 2424
rect 17770 2388 17800 2424
rect 17914 2388 17944 2424
rect 18058 2388 18088 2424
rect 18202 2388 18232 2424
rect 18346 2388 18376 2424
rect 18490 2388 18520 2424
rect 18634 2388 18664 2424
rect 18778 2388 18808 2424
rect 18922 2388 18952 2424
rect 19066 2388 19096 2424
rect 19210 2388 19240 2424
rect 19354 2388 19384 2424
rect 19498 2388 19528 2424
rect 19642 2388 19672 2424
rect 19786 2388 19816 2424
rect 19930 2388 19960 2424
rect 776 1608 806 1644
rect 920 1608 950 1644
rect 1352 1608 1382 1644
rect 1496 1608 1526 1644
rect 1928 1608 1958 1644
rect 2072 1608 2102 1644
rect 3080 1608 3110 1644
rect 3224 1608 3254 1644
rect 3656 1608 3686 1644
rect 3800 1608 3830 1644
rect 4232 1608 4262 1644
rect 4376 1608 4406 1644
rect 5960 1608 5990 1644
rect 6104 1608 6134 1644
rect 6536 1608 6566 1644
rect 6680 1608 6710 1644
rect 7112 1608 7142 1644
rect 7256 1608 7286 1644
rect 7688 1608 7718 1644
rect 7832 1608 7862 1644
rect 8264 1608 8294 1644
rect 8408 1608 8438 1644
rect 9416 1608 9446 1644
rect 9560 1608 9590 1644
rect 9992 1608 10022 1644
rect 10136 1608 10166 1644
rect 10568 1608 10598 1644
rect 10712 1608 10742 1644
rect 11144 1608 11174 1644
rect 11288 1608 11318 1644
rect 12008 1608 12038 1644
rect 12152 1608 12182 1644
rect 12584 1608 12614 1644
rect 12728 1608 12758 1644
rect 13160 1608 13190 1644
rect 13304 1608 13334 1644
rect 13736 1608 13766 1644
rect 13880 1608 13910 1644
rect 14888 1608 14918 1644
rect 15032 1608 15062 1644
rect 15466 1608 15496 1644
rect 15610 1608 15640 1644
rect 16040 1608 16070 1644
rect 16184 1608 16214 1644
rect 16328 1608 16358 1644
rect 16472 1608 16502 1644
rect 17480 1608 17510 1644
rect 17624 1608 17654 1644
rect 17768 1608 17798 1644
rect 17912 1608 17942 1644
rect 18056 1608 18086 1644
rect 18200 1608 18230 1644
rect 18344 1608 18374 1644
rect 18488 1608 18518 1644
rect 18632 1608 18662 1644
rect 18776 1608 18806 1644
rect 18920 1608 18950 1644
rect 19064 1608 19094 1644
rect 19208 1608 19238 1644
rect 19352 1608 19382 1644
rect 19496 1608 19526 1644
rect 19640 1608 19670 1644
rect 19784 1608 19814 1644
rect 19928 1608 19958 1644
rect 20072 1608 20102 1644
rect 20216 1608 20246 1644
rect 20360 1608 20390 1644
rect 20504 1608 20534 1644
rect 20648 1608 20678 1644
rect 20792 1608 20822 1644
rect 776 1332 806 1368
rect 920 1332 950 1368
rect 776 1313 950 1332
rect 776 1279 796 1313
rect 830 1279 904 1313
rect 938 1279 950 1313
rect 776 1260 950 1279
rect 1352 1332 1382 1368
rect 1496 1332 1526 1368
rect 1352 1313 1526 1332
rect 1352 1279 1372 1313
rect 1406 1279 1480 1313
rect 1514 1279 1526 1313
rect 1352 1260 1526 1279
rect 1928 1332 1958 1368
rect 2072 1332 2102 1368
rect 1928 1313 2102 1332
rect 1928 1279 1948 1313
rect 1982 1279 2056 1313
rect 2090 1279 2102 1313
rect 1928 1260 2102 1279
rect 3080 1332 3110 1368
rect 3224 1332 3254 1368
rect 3080 1313 3254 1332
rect 3080 1279 3100 1313
rect 3134 1279 3208 1313
rect 3242 1279 3254 1313
rect 3080 1260 3254 1279
rect 3656 1332 3686 1368
rect 3800 1332 3830 1368
rect 3656 1313 3830 1332
rect 3656 1279 3676 1313
rect 3710 1279 3784 1313
rect 3818 1279 3830 1313
rect 3656 1260 3830 1279
rect 4232 1332 4262 1368
rect 4376 1332 4406 1368
rect 4232 1313 4406 1332
rect 4232 1279 4252 1313
rect 4286 1279 4360 1313
rect 4394 1279 4406 1313
rect 4232 1260 4406 1279
rect 5960 1332 5990 1368
rect 6104 1332 6134 1368
rect 5960 1313 6134 1332
rect 5960 1279 5980 1313
rect 6014 1279 6088 1313
rect 6122 1279 6134 1313
rect 5960 1260 6134 1279
rect 6536 1332 6566 1368
rect 6680 1332 6710 1368
rect 6536 1313 6710 1332
rect 6536 1279 6556 1313
rect 6590 1279 6664 1313
rect 6698 1279 6710 1313
rect 6536 1260 6710 1279
rect 7112 1332 7142 1368
rect 7256 1332 7286 1368
rect 7112 1313 7286 1332
rect 7112 1279 7132 1313
rect 7166 1279 7240 1313
rect 7274 1279 7286 1313
rect 7112 1260 7286 1279
rect 7688 1332 7718 1368
rect 7832 1332 7862 1368
rect 8264 1332 8294 1368
rect 7688 1313 7862 1332
rect 7688 1279 7708 1313
rect 7742 1279 7816 1313
rect 7850 1279 7862 1313
rect 7688 1260 7862 1279
rect 8174 1314 8294 1332
rect 8174 1278 8196 1314
rect 8232 1278 8294 1314
rect 8174 1260 8294 1278
rect 8408 1332 8438 1368
rect 9416 1332 9446 1368
rect 9560 1332 9590 1368
rect 8408 1314 8528 1332
rect 8408 1278 8474 1314
rect 8510 1278 8528 1314
rect 8408 1260 8528 1278
rect 9416 1313 9590 1332
rect 9416 1279 9436 1313
rect 9470 1279 9544 1313
rect 9578 1279 9590 1313
rect 9416 1260 9590 1279
rect 9992 1332 10022 1368
rect 10136 1332 10166 1368
rect 9992 1313 10166 1332
rect 9992 1279 10012 1313
rect 10046 1279 10120 1313
rect 10154 1279 10166 1313
rect 9992 1260 10166 1279
rect 10568 1332 10598 1368
rect 10712 1332 10742 1368
rect 11144 1332 11174 1368
rect 10568 1313 10742 1332
rect 10568 1279 10588 1313
rect 10622 1279 10696 1313
rect 10730 1279 10742 1313
rect 10568 1260 10742 1279
rect 11054 1314 11174 1332
rect 11054 1278 11076 1314
rect 11112 1278 11174 1314
rect 11054 1260 11174 1278
rect 11288 1332 11318 1368
rect 12008 1332 12038 1368
rect 12152 1332 12182 1368
rect 11288 1314 11408 1332
rect 11288 1278 11354 1314
rect 11390 1278 11408 1314
rect 11288 1260 11408 1278
rect 12008 1313 12182 1332
rect 12008 1279 12028 1313
rect 12062 1279 12136 1313
rect 12170 1279 12182 1313
rect 12008 1260 12182 1279
rect 12584 1332 12614 1368
rect 12728 1332 12758 1368
rect 12584 1313 12758 1332
rect 12584 1279 12604 1313
rect 12638 1279 12712 1313
rect 12746 1279 12758 1313
rect 12584 1260 12758 1279
rect 13160 1332 13190 1368
rect 13304 1332 13334 1368
rect 13160 1313 13334 1332
rect 13160 1279 13180 1313
rect 13214 1279 13288 1313
rect 13322 1279 13334 1313
rect 13160 1260 13334 1279
rect 13736 1332 13766 1368
rect 13880 1332 13910 1368
rect 13736 1313 13910 1332
rect 13736 1279 13756 1313
rect 13790 1279 13864 1313
rect 13898 1279 13910 1313
rect 13736 1260 13910 1279
rect 14888 1332 14918 1368
rect 15032 1332 15062 1368
rect 14888 1313 15062 1332
rect 14888 1279 14908 1313
rect 14942 1279 15016 1313
rect 15050 1279 15062 1313
rect 14888 1260 15062 1279
rect 15466 1332 15496 1368
rect 15610 1332 15640 1368
rect 15466 1313 15640 1332
rect 15466 1279 15478 1313
rect 15512 1279 15586 1313
rect 15620 1279 15640 1313
rect 15466 1260 15640 1279
rect 16040 1332 16070 1368
rect 16184 1332 16214 1368
rect 16040 1313 16214 1332
rect 16040 1279 16060 1313
rect 16094 1279 16168 1313
rect 16202 1279 16214 1313
rect 16040 1260 16214 1279
rect 16328 1332 16358 1368
rect 16472 1332 16502 1368
rect 16328 1313 16502 1332
rect 16328 1279 16348 1313
rect 16382 1279 16456 1313
rect 16490 1279 16502 1313
rect 16328 1260 16502 1279
rect 17480 1332 17510 1368
rect 17624 1332 17654 1368
rect 17480 1313 17654 1332
rect 17480 1279 17500 1313
rect 17534 1279 17608 1313
rect 17642 1279 17654 1313
rect 17480 1260 17654 1279
rect 17768 1332 17798 1368
rect 17912 1332 17942 1368
rect 17768 1313 17942 1332
rect 17768 1279 17788 1313
rect 17822 1279 17896 1313
rect 17930 1279 17942 1313
rect 17768 1260 17942 1279
rect 18056 1332 18086 1368
rect 18200 1332 18230 1368
rect 18056 1313 18230 1332
rect 18056 1279 18076 1313
rect 18110 1279 18184 1313
rect 18218 1279 18230 1313
rect 18056 1260 18230 1279
rect 18344 1332 18374 1368
rect 18488 1332 18518 1368
rect 18344 1313 18518 1332
rect 18344 1279 18364 1313
rect 18398 1279 18472 1313
rect 18506 1279 18518 1313
rect 18344 1260 18518 1279
rect 18632 1332 18662 1368
rect 18776 1332 18806 1368
rect 18632 1313 18806 1332
rect 18632 1279 18652 1313
rect 18686 1279 18760 1313
rect 18794 1279 18806 1313
rect 18632 1260 18806 1279
rect 18920 1332 18950 1368
rect 19064 1332 19094 1368
rect 18920 1313 19094 1332
rect 18920 1279 18940 1313
rect 18974 1279 19048 1313
rect 19082 1279 19094 1313
rect 18920 1260 19094 1279
rect 19208 1332 19238 1368
rect 19352 1332 19382 1368
rect 19208 1313 19382 1332
rect 19208 1279 19228 1313
rect 19262 1279 19336 1313
rect 19370 1279 19382 1313
rect 19208 1260 19382 1279
rect 19496 1332 19526 1368
rect 19640 1332 19670 1368
rect 19496 1313 19670 1332
rect 19496 1279 19516 1313
rect 19550 1279 19624 1313
rect 19658 1279 19670 1313
rect 19496 1260 19670 1279
rect 19784 1332 19814 1368
rect 19928 1332 19958 1368
rect 19784 1313 19958 1332
rect 19784 1279 19804 1313
rect 19838 1279 19912 1313
rect 19946 1279 19958 1313
rect 19784 1260 19958 1279
rect 20072 1332 20102 1368
rect 20216 1332 20246 1368
rect 20072 1313 20246 1332
rect 20072 1279 20092 1313
rect 20126 1279 20200 1313
rect 20234 1279 20246 1313
rect 20072 1260 20246 1279
rect 20360 1332 20390 1368
rect 20504 1332 20534 1368
rect 20360 1313 20534 1332
rect 20360 1279 20380 1313
rect 20414 1279 20488 1313
rect 20522 1279 20534 1313
rect 20360 1260 20534 1279
rect 20648 1332 20678 1368
rect 20792 1332 20822 1368
rect 20648 1313 20822 1332
rect 20648 1279 20668 1313
rect 20702 1279 20776 1313
rect 20810 1279 20822 1313
rect 20648 1260 20822 1279
rect 776 737 950 756
rect 776 703 796 737
rect 830 703 904 737
rect 938 703 950 737
rect 776 684 950 703
rect 776 648 806 684
rect 920 648 950 684
rect 1352 737 1526 756
rect 1352 703 1372 737
rect 1406 703 1480 737
rect 1514 703 1526 737
rect 1352 684 1526 703
rect 1352 648 1382 684
rect 1496 648 1526 684
rect 1928 737 2102 756
rect 1928 703 1948 737
rect 1982 703 2056 737
rect 2090 703 2102 737
rect 1928 684 2102 703
rect 1928 648 1958 684
rect 2072 648 2102 684
rect 3080 737 3254 756
rect 3080 703 3100 737
rect 3134 703 3208 737
rect 3242 703 3254 737
rect 3080 684 3254 703
rect 3080 648 3110 684
rect 3224 648 3254 684
rect 3656 737 3830 756
rect 3656 703 3676 737
rect 3710 703 3784 737
rect 3818 703 3830 737
rect 3656 684 3830 703
rect 3656 648 3686 684
rect 3800 648 3830 684
rect 4232 737 4406 756
rect 4232 703 4252 737
rect 4286 703 4360 737
rect 4394 703 4406 737
rect 4232 684 4406 703
rect 4232 648 4262 684
rect 4376 648 4406 684
rect 5960 737 6134 756
rect 5960 703 5980 737
rect 6014 703 6088 737
rect 6122 703 6134 737
rect 5960 684 6134 703
rect 5960 648 5990 684
rect 6104 648 6134 684
rect 6536 737 6710 756
rect 6536 703 6556 737
rect 6590 703 6664 737
rect 6698 703 6710 737
rect 6536 684 6710 703
rect 6536 648 6566 684
rect 6680 648 6710 684
rect 7112 737 7286 756
rect 7112 703 7132 737
rect 7166 703 7240 737
rect 7274 703 7286 737
rect 7112 684 7286 703
rect 7112 648 7142 684
rect 7256 648 7286 684
rect 7688 737 7862 756
rect 7688 703 7708 737
rect 7742 703 7816 737
rect 7850 703 7862 737
rect 7688 684 7862 703
rect 8174 738 8294 756
rect 8174 702 8196 738
rect 8232 702 8294 738
rect 8174 684 8294 702
rect 7688 648 7718 684
rect 7832 648 7862 684
rect 8264 648 8294 684
rect 8408 738 8528 756
rect 8408 702 8480 738
rect 8516 702 8528 738
rect 8408 684 8528 702
rect 9416 737 9590 756
rect 9416 703 9436 737
rect 9470 703 9544 737
rect 9578 703 9590 737
rect 9416 684 9590 703
rect 8408 648 8438 684
rect 9416 648 9446 684
rect 9560 648 9590 684
rect 9992 737 10166 756
rect 9992 703 10012 737
rect 10046 703 10120 737
rect 10154 703 10166 737
rect 9992 684 10166 703
rect 9992 648 10022 684
rect 10136 648 10166 684
rect 10568 737 10742 756
rect 10568 703 10588 737
rect 10622 703 10696 737
rect 10730 703 10742 737
rect 10568 684 10742 703
rect 11054 738 11174 756
rect 11054 702 11076 738
rect 11112 702 11174 738
rect 11054 684 11174 702
rect 10568 648 10598 684
rect 10712 648 10742 684
rect 11144 648 11174 684
rect 11288 738 11408 756
rect 11288 702 11360 738
rect 11396 702 11408 738
rect 11288 684 11408 702
rect 12008 737 12182 756
rect 12008 703 12028 737
rect 12062 703 12136 737
rect 12170 703 12182 737
rect 12008 684 12182 703
rect 11288 648 11318 684
rect 12008 648 12038 684
rect 12152 648 12182 684
rect 12584 737 12758 756
rect 12584 703 12604 737
rect 12638 703 12712 737
rect 12746 703 12758 737
rect 12584 684 12758 703
rect 12584 648 12614 684
rect 12728 648 12758 684
rect 13160 737 13334 756
rect 13160 703 13180 737
rect 13214 703 13288 737
rect 13322 703 13334 737
rect 13160 684 13334 703
rect 13160 648 13190 684
rect 13304 648 13334 684
rect 13736 737 13910 756
rect 13736 703 13756 737
rect 13790 703 13864 737
rect 13898 703 13910 737
rect 13736 684 13910 703
rect 13736 648 13766 684
rect 13880 648 13910 684
rect 14888 737 15062 756
rect 14888 703 14908 737
rect 14942 703 15016 737
rect 15050 703 15062 737
rect 14888 684 15062 703
rect 14888 648 14918 684
rect 15032 648 15062 684
rect 15466 737 15640 756
rect 15466 703 15478 737
rect 15512 703 15586 737
rect 15620 703 15640 737
rect 15466 684 15640 703
rect 15466 648 15496 684
rect 15610 648 15640 684
rect 16040 737 16214 756
rect 16040 703 16060 737
rect 16094 703 16168 737
rect 16202 703 16214 737
rect 16040 684 16214 703
rect 16040 648 16070 684
rect 16184 648 16214 684
rect 16328 737 16502 756
rect 16328 703 16348 737
rect 16382 703 16456 737
rect 16490 703 16502 737
rect 16328 684 16502 703
rect 16328 648 16358 684
rect 16472 648 16502 684
rect 17480 737 17654 756
rect 17480 703 17500 737
rect 17534 703 17608 737
rect 17642 703 17654 737
rect 17480 684 17654 703
rect 17480 648 17510 684
rect 17624 648 17654 684
rect 17768 737 17942 756
rect 17768 703 17788 737
rect 17822 703 17896 737
rect 17930 703 17942 737
rect 17768 684 17942 703
rect 17768 648 17798 684
rect 17912 648 17942 684
rect 18056 737 18230 756
rect 18056 703 18076 737
rect 18110 703 18184 737
rect 18218 703 18230 737
rect 18056 684 18230 703
rect 18056 648 18086 684
rect 18200 648 18230 684
rect 18344 737 18518 756
rect 18344 703 18364 737
rect 18398 703 18472 737
rect 18506 703 18518 737
rect 18344 684 18518 703
rect 18344 648 18374 684
rect 18488 648 18518 684
rect 18632 737 18806 756
rect 18632 703 18652 737
rect 18686 703 18760 737
rect 18794 703 18806 737
rect 18632 684 18806 703
rect 18632 648 18662 684
rect 18776 648 18806 684
rect 18920 737 19094 756
rect 18920 703 18940 737
rect 18974 703 19048 737
rect 19082 703 19094 737
rect 18920 684 19094 703
rect 18920 648 18950 684
rect 19064 648 19094 684
rect 19208 737 19382 756
rect 19208 703 19228 737
rect 19262 703 19336 737
rect 19370 703 19382 737
rect 19208 684 19382 703
rect 19208 648 19238 684
rect 19352 648 19382 684
rect 19496 737 19670 756
rect 19496 703 19516 737
rect 19550 703 19624 737
rect 19658 703 19670 737
rect 19496 684 19670 703
rect 19496 648 19526 684
rect 19640 648 19670 684
rect 19784 737 19958 756
rect 19784 703 19804 737
rect 19838 703 19912 737
rect 19946 703 19958 737
rect 19784 684 19958 703
rect 19784 648 19814 684
rect 19928 648 19958 684
rect 20072 737 20246 756
rect 20072 703 20092 737
rect 20126 703 20200 737
rect 20234 703 20246 737
rect 20072 684 20246 703
rect 20072 648 20102 684
rect 20216 648 20246 684
rect 20360 737 20534 756
rect 20360 703 20380 737
rect 20414 703 20488 737
rect 20522 703 20534 737
rect 20360 684 20534 703
rect 20360 648 20390 684
rect 20504 648 20534 684
rect 20648 737 20822 756
rect 20648 703 20668 737
rect 20702 703 20776 737
rect 20810 703 20822 737
rect 20648 684 20822 703
rect 20648 648 20678 684
rect 20792 648 20822 684
rect 776 132 806 168
rect 920 132 950 168
rect 1352 132 1382 168
rect 1496 132 1526 168
rect 1928 132 1958 168
rect 2072 132 2102 168
rect 3080 132 3110 168
rect 3224 132 3254 168
rect 3656 132 3686 168
rect 3800 132 3830 168
rect 4232 132 4262 168
rect 4376 132 4406 168
rect 5960 132 5990 168
rect 6104 132 6134 168
rect 6536 132 6566 168
rect 6680 132 6710 168
rect 7112 132 7142 168
rect 7256 132 7286 168
rect 7688 132 7718 168
rect 7832 132 7862 168
rect 8264 132 8294 168
rect 8408 132 8438 168
rect 9416 132 9446 168
rect 9560 132 9590 168
rect 9992 132 10022 168
rect 10136 132 10166 168
rect 10568 132 10598 168
rect 10712 132 10742 168
rect 11144 132 11174 168
rect 11288 132 11318 168
rect 12008 132 12038 168
rect 12152 132 12182 168
rect 12584 132 12614 168
rect 12728 132 12758 168
rect 13160 132 13190 168
rect 13304 132 13334 168
rect 13736 132 13766 168
rect 13880 132 13910 168
rect 14888 132 14918 168
rect 15032 132 15062 168
rect 15466 132 15496 168
rect 15610 132 15640 168
rect 16040 132 16070 168
rect 16184 132 16214 168
rect 16328 132 16358 168
rect 16472 132 16502 168
rect 17480 132 17510 168
rect 17624 132 17654 168
rect 17768 132 17798 168
rect 17912 132 17942 168
rect 18056 132 18086 168
rect 18200 132 18230 168
rect 18344 132 18374 168
rect 18488 132 18518 168
rect 18632 132 18662 168
rect 18776 132 18806 168
rect 18920 132 18950 168
rect 19064 132 19094 168
rect 19208 132 19238 168
rect 19352 132 19382 168
rect 19496 132 19526 168
rect 19640 132 19670 168
rect 19784 132 19814 168
rect 19928 132 19958 168
rect 20072 132 20102 168
rect 20216 132 20246 168
rect 20360 132 20390 168
rect 20504 132 20534 168
rect 20648 132 20678 168
rect 20792 132 20822 168
<< polycont >>
rect 790 3295 824 3329
rect 898 3295 932 3329
rect 1366 3295 1400 3329
rect 1474 3295 1508 3329
rect 1942 3295 1976 3329
rect 2050 3295 2084 3329
rect 2518 3295 2552 3329
rect 2626 3295 2660 3329
rect 3100 3295 3134 3329
rect 3208 3295 3242 3329
rect 4252 3295 4286 3329
rect 4360 3295 4394 3329
rect 4828 3295 4862 3329
rect 4936 3295 4970 3329
rect 5404 3295 5438 3329
rect 5512 3295 5546 3329
rect 5980 3295 6014 3329
rect 6088 3295 6122 3329
rect 6468 3294 6504 3330
rect 6752 3294 6788 3330
rect 7708 3295 7742 3329
rect 7816 3295 7850 3329
rect 8284 3295 8318 3329
rect 8392 3295 8426 3329
rect 8860 3295 8894 3329
rect 8968 3295 9002 3329
rect 9348 3294 9384 3330
rect 9632 3294 9668 3330
rect 10300 3295 10334 3329
rect 10408 3295 10442 3329
rect 10876 3295 10910 3329
rect 10984 3295 11018 3329
rect 12028 3295 12062 3329
rect 12136 3295 12170 3329
rect 12604 3295 12638 3329
rect 12712 3295 12746 3329
rect 13756 3295 13790 3329
rect 13864 3295 13898 3329
rect 14332 3295 14366 3329
rect 14440 3295 14474 3329
rect 14908 3295 14942 3329
rect 15016 3295 15050 3329
rect 16630 3295 16664 3329
rect 16738 3295 16772 3329
rect 16918 3295 16952 3329
rect 17026 3295 17060 3329
rect 17206 3295 17240 3329
rect 17314 3295 17348 3329
rect 17494 3295 17528 3329
rect 17602 3295 17636 3329
rect 17782 3295 17816 3329
rect 17890 3295 17924 3329
rect 18070 3295 18104 3329
rect 18178 3295 18212 3329
rect 18358 3295 18392 3329
rect 18466 3295 18500 3329
rect 18646 3295 18680 3329
rect 18754 3295 18788 3329
rect 18934 3295 18968 3329
rect 19042 3295 19076 3329
rect 19222 3295 19256 3329
rect 19330 3295 19364 3329
rect 19510 3295 19544 3329
rect 19618 3295 19652 3329
rect 19798 3295 19832 3329
rect 19906 3295 19940 3329
rect 790 2719 824 2753
rect 898 2719 932 2753
rect 1366 2719 1400 2753
rect 1474 2719 1508 2753
rect 1942 2719 1976 2753
rect 2050 2719 2084 2753
rect 2518 2719 2552 2753
rect 2626 2719 2660 2753
rect 3100 2719 3134 2753
rect 3208 2719 3242 2753
rect 4252 2719 4286 2753
rect 4360 2719 4394 2753
rect 4828 2719 4862 2753
rect 4936 2719 4970 2753
rect 5404 2719 5438 2753
rect 5512 2719 5546 2753
rect 5980 2719 6014 2753
rect 6088 2719 6122 2753
rect 6468 2718 6504 2754
rect 6746 2718 6782 2754
rect 7708 2719 7742 2753
rect 7816 2719 7850 2753
rect 8284 2719 8318 2753
rect 8392 2719 8426 2753
rect 8860 2719 8894 2753
rect 8968 2719 9002 2753
rect 9348 2718 9384 2754
rect 9626 2718 9662 2754
rect 10300 2719 10334 2753
rect 10408 2719 10442 2753
rect 10876 2719 10910 2753
rect 10984 2719 11018 2753
rect 12028 2719 12062 2753
rect 12136 2719 12170 2753
rect 12604 2719 12638 2753
rect 12712 2719 12746 2753
rect 13756 2719 13790 2753
rect 13864 2719 13898 2753
rect 14332 2719 14366 2753
rect 14440 2719 14474 2753
rect 14908 2719 14942 2753
rect 15016 2719 15050 2753
rect 16630 2719 16664 2753
rect 16738 2719 16772 2753
rect 16918 2719 16952 2753
rect 17026 2719 17060 2753
rect 17206 2719 17240 2753
rect 17314 2719 17348 2753
rect 17494 2719 17528 2753
rect 17602 2719 17636 2753
rect 17782 2719 17816 2753
rect 17890 2719 17924 2753
rect 18070 2719 18104 2753
rect 18178 2719 18212 2753
rect 18358 2719 18392 2753
rect 18466 2719 18500 2753
rect 18646 2719 18680 2753
rect 18754 2719 18788 2753
rect 18934 2719 18968 2753
rect 19042 2719 19076 2753
rect 19222 2719 19256 2753
rect 19330 2719 19364 2753
rect 19510 2719 19544 2753
rect 19618 2719 19652 2753
rect 19798 2719 19832 2753
rect 19906 2719 19940 2753
rect 796 1279 830 1313
rect 904 1279 938 1313
rect 1372 1279 1406 1313
rect 1480 1279 1514 1313
rect 1948 1279 1982 1313
rect 2056 1279 2090 1313
rect 3100 1279 3134 1313
rect 3208 1279 3242 1313
rect 3676 1279 3710 1313
rect 3784 1279 3818 1313
rect 4252 1279 4286 1313
rect 4360 1279 4394 1313
rect 5980 1279 6014 1313
rect 6088 1279 6122 1313
rect 6556 1279 6590 1313
rect 6664 1279 6698 1313
rect 7132 1279 7166 1313
rect 7240 1279 7274 1313
rect 7708 1279 7742 1313
rect 7816 1279 7850 1313
rect 8196 1278 8232 1314
rect 8474 1278 8510 1314
rect 9436 1279 9470 1313
rect 9544 1279 9578 1313
rect 10012 1279 10046 1313
rect 10120 1279 10154 1313
rect 10588 1279 10622 1313
rect 10696 1279 10730 1313
rect 11076 1278 11112 1314
rect 11354 1278 11390 1314
rect 12028 1279 12062 1313
rect 12136 1279 12170 1313
rect 12604 1279 12638 1313
rect 12712 1279 12746 1313
rect 13180 1279 13214 1313
rect 13288 1279 13322 1313
rect 13756 1279 13790 1313
rect 13864 1279 13898 1313
rect 14908 1279 14942 1313
rect 15016 1279 15050 1313
rect 15478 1279 15512 1313
rect 15586 1279 15620 1313
rect 16060 1279 16094 1313
rect 16168 1279 16202 1313
rect 16348 1279 16382 1313
rect 16456 1279 16490 1313
rect 17500 1279 17534 1313
rect 17608 1279 17642 1313
rect 17788 1279 17822 1313
rect 17896 1279 17930 1313
rect 18076 1279 18110 1313
rect 18184 1279 18218 1313
rect 18364 1279 18398 1313
rect 18472 1279 18506 1313
rect 18652 1279 18686 1313
rect 18760 1279 18794 1313
rect 18940 1279 18974 1313
rect 19048 1279 19082 1313
rect 19228 1279 19262 1313
rect 19336 1279 19370 1313
rect 19516 1279 19550 1313
rect 19624 1279 19658 1313
rect 19804 1279 19838 1313
rect 19912 1279 19946 1313
rect 20092 1279 20126 1313
rect 20200 1279 20234 1313
rect 20380 1279 20414 1313
rect 20488 1279 20522 1313
rect 20668 1279 20702 1313
rect 20776 1279 20810 1313
rect 796 703 830 737
rect 904 703 938 737
rect 1372 703 1406 737
rect 1480 703 1514 737
rect 1948 703 1982 737
rect 2056 703 2090 737
rect 3100 703 3134 737
rect 3208 703 3242 737
rect 3676 703 3710 737
rect 3784 703 3818 737
rect 4252 703 4286 737
rect 4360 703 4394 737
rect 5980 703 6014 737
rect 6088 703 6122 737
rect 6556 703 6590 737
rect 6664 703 6698 737
rect 7132 703 7166 737
rect 7240 703 7274 737
rect 7708 703 7742 737
rect 7816 703 7850 737
rect 8196 702 8232 738
rect 8480 702 8516 738
rect 9436 703 9470 737
rect 9544 703 9578 737
rect 10012 703 10046 737
rect 10120 703 10154 737
rect 10588 703 10622 737
rect 10696 703 10730 737
rect 11076 702 11112 738
rect 11360 702 11396 738
rect 12028 703 12062 737
rect 12136 703 12170 737
rect 12604 703 12638 737
rect 12712 703 12746 737
rect 13180 703 13214 737
rect 13288 703 13322 737
rect 13756 703 13790 737
rect 13864 703 13898 737
rect 14908 703 14942 737
rect 15016 703 15050 737
rect 15478 703 15512 737
rect 15586 703 15620 737
rect 16060 703 16094 737
rect 16168 703 16202 737
rect 16348 703 16382 737
rect 16456 703 16490 737
rect 17500 703 17534 737
rect 17608 703 17642 737
rect 17788 703 17822 737
rect 17896 703 17930 737
rect 18076 703 18110 737
rect 18184 703 18218 737
rect 18364 703 18398 737
rect 18472 703 18506 737
rect 18652 703 18686 737
rect 18760 703 18794 737
rect 18940 703 18974 737
rect 19048 703 19082 737
rect 19228 703 19262 737
rect 19336 703 19370 737
rect 19516 703 19550 737
rect 19624 703 19658 737
rect 19804 703 19838 737
rect 19912 703 19946 737
rect 20092 703 20126 737
rect 20200 703 20234 737
rect 20380 703 20414 737
rect 20488 703 20522 737
rect 20668 703 20702 737
rect 20776 703 20810 737
<< locali >>
rect 690 3794 750 3810
rect 690 3754 700 3794
rect 740 3754 750 3794
rect 114 3704 174 3728
rect 114 3552 124 3704
rect 164 3552 174 3704
rect 114 3528 174 3552
rect 258 3704 318 3728
rect 258 3552 268 3704
rect 308 3552 318 3704
rect 258 3528 318 3552
rect 402 3704 462 3728
rect 402 3552 412 3704
rect 452 3552 462 3704
rect 402 3528 462 3552
rect 690 3694 750 3754
rect 690 3654 700 3694
rect 740 3654 750 3694
rect 690 3594 750 3654
rect 690 3554 700 3594
rect 740 3554 750 3594
rect 690 3494 750 3554
rect 690 3454 700 3494
rect 740 3454 750 3494
rect 690 3438 750 3454
rect 834 3794 894 3810
rect 834 3754 844 3794
rect 884 3754 894 3794
rect 834 3694 894 3754
rect 834 3654 844 3694
rect 884 3654 894 3694
rect 834 3594 894 3654
rect 834 3554 844 3594
rect 884 3554 894 3594
rect 834 3494 894 3554
rect 834 3454 844 3494
rect 884 3454 894 3494
rect 834 3438 894 3454
rect 978 3794 1038 3810
rect 978 3754 988 3794
rect 1028 3754 1038 3794
rect 978 3694 1038 3754
rect 978 3654 988 3694
rect 1028 3654 1038 3694
rect 978 3594 1038 3654
rect 978 3554 988 3594
rect 1028 3554 1038 3594
rect 978 3494 1038 3554
rect 978 3454 988 3494
rect 1028 3454 1038 3494
rect 978 3438 1038 3454
rect 1266 3794 1326 3810
rect 1266 3754 1276 3794
rect 1316 3754 1326 3794
rect 1266 3694 1326 3754
rect 1266 3654 1276 3694
rect 1316 3654 1326 3694
rect 1266 3594 1326 3654
rect 1266 3554 1276 3594
rect 1316 3554 1326 3594
rect 1266 3494 1326 3554
rect 1266 3454 1276 3494
rect 1316 3454 1326 3494
rect 1266 3438 1326 3454
rect 1410 3794 1470 3810
rect 1410 3754 1420 3794
rect 1460 3754 1470 3794
rect 1410 3694 1470 3754
rect 1410 3654 1420 3694
rect 1460 3654 1470 3694
rect 1410 3594 1470 3654
rect 1410 3554 1420 3594
rect 1460 3554 1470 3594
rect 1410 3494 1470 3554
rect 1410 3454 1420 3494
rect 1460 3454 1470 3494
rect 1410 3438 1470 3454
rect 1554 3794 1614 3810
rect 1554 3754 1564 3794
rect 1604 3754 1614 3794
rect 1554 3694 1614 3754
rect 1554 3654 1564 3694
rect 1604 3654 1614 3694
rect 1554 3594 1614 3654
rect 1554 3554 1564 3594
rect 1604 3554 1614 3594
rect 1554 3494 1614 3554
rect 1554 3454 1564 3494
rect 1604 3454 1614 3494
rect 1554 3438 1614 3454
rect 1842 3794 1902 3810
rect 1842 3754 1852 3794
rect 1892 3754 1902 3794
rect 1842 3694 1902 3754
rect 1842 3654 1852 3694
rect 1892 3654 1902 3694
rect 1842 3594 1902 3654
rect 1842 3554 1852 3594
rect 1892 3554 1902 3594
rect 1842 3494 1902 3554
rect 1842 3454 1852 3494
rect 1892 3454 1902 3494
rect 1842 3438 1902 3454
rect 1986 3794 2046 3810
rect 1986 3754 1996 3794
rect 2036 3754 2046 3794
rect 1986 3694 2046 3754
rect 1986 3654 1996 3694
rect 2036 3654 2046 3694
rect 1986 3594 2046 3654
rect 1986 3554 1996 3594
rect 2036 3554 2046 3594
rect 1986 3494 2046 3554
rect 1986 3454 1996 3494
rect 2036 3454 2046 3494
rect 1986 3438 2046 3454
rect 2130 3794 2190 3810
rect 2130 3754 2140 3794
rect 2180 3754 2190 3794
rect 2130 3694 2190 3754
rect 2130 3654 2140 3694
rect 2180 3654 2190 3694
rect 2130 3594 2190 3654
rect 2130 3554 2140 3594
rect 2180 3554 2190 3594
rect 2130 3494 2190 3554
rect 2130 3454 2140 3494
rect 2180 3454 2190 3494
rect 2130 3438 2190 3454
rect 2418 3794 2478 3810
rect 2418 3754 2428 3794
rect 2468 3754 2478 3794
rect 2418 3694 2478 3754
rect 2418 3654 2428 3694
rect 2468 3654 2478 3694
rect 2418 3594 2478 3654
rect 2418 3554 2428 3594
rect 2468 3554 2478 3594
rect 2418 3494 2478 3554
rect 2418 3454 2428 3494
rect 2468 3454 2478 3494
rect 2418 3438 2478 3454
rect 2562 3794 2622 3810
rect 2562 3754 2572 3794
rect 2612 3754 2622 3794
rect 2562 3694 2622 3754
rect 2562 3654 2572 3694
rect 2612 3654 2622 3694
rect 2562 3594 2622 3654
rect 2562 3554 2572 3594
rect 2612 3554 2622 3594
rect 2562 3494 2622 3554
rect 2562 3454 2572 3494
rect 2612 3454 2622 3494
rect 2562 3438 2622 3454
rect 2706 3794 2766 3810
rect 2706 3754 2716 3794
rect 2756 3754 2766 3794
rect 2706 3694 2766 3754
rect 2706 3654 2716 3694
rect 2756 3654 2766 3694
rect 2706 3594 2766 3654
rect 2706 3554 2716 3594
rect 2756 3554 2766 3594
rect 2706 3494 2766 3554
rect 2706 3454 2716 3494
rect 2756 3454 2766 3494
rect 2706 3438 2766 3454
rect 2994 3794 3054 3810
rect 2994 3754 3004 3794
rect 3044 3754 3054 3794
rect 2994 3694 3054 3754
rect 2994 3654 3004 3694
rect 3044 3654 3054 3694
rect 2994 3594 3054 3654
rect 2994 3554 3004 3594
rect 3044 3554 3054 3594
rect 2994 3494 3054 3554
rect 2994 3454 3004 3494
rect 3044 3454 3054 3494
rect 2994 3438 3054 3454
rect 3138 3794 3198 3810
rect 3138 3754 3148 3794
rect 3188 3754 3198 3794
rect 3138 3694 3198 3754
rect 3138 3654 3148 3694
rect 3188 3654 3198 3694
rect 3138 3594 3198 3654
rect 3138 3554 3148 3594
rect 3188 3554 3198 3594
rect 3138 3494 3198 3554
rect 3138 3454 3148 3494
rect 3188 3454 3198 3494
rect 3138 3438 3198 3454
rect 3282 3794 3342 3810
rect 3282 3754 3292 3794
rect 3332 3754 3342 3794
rect 3282 3694 3342 3754
rect 4146 3794 4206 3810
rect 4146 3754 4156 3794
rect 4196 3754 4206 3794
rect 3282 3654 3292 3694
rect 3332 3654 3342 3694
rect 3282 3594 3342 3654
rect 3282 3554 3292 3594
rect 3332 3554 3342 3594
rect 3282 3494 3342 3554
rect 3570 3704 3630 3728
rect 3570 3552 3580 3704
rect 3620 3552 3630 3704
rect 3570 3528 3630 3552
rect 3714 3704 3774 3728
rect 3714 3552 3724 3704
rect 3764 3552 3774 3704
rect 3714 3528 3774 3552
rect 3858 3704 3918 3728
rect 3858 3552 3868 3704
rect 3908 3552 3918 3704
rect 3858 3528 3918 3552
rect 4146 3694 4206 3754
rect 4146 3654 4156 3694
rect 4196 3654 4206 3694
rect 4146 3594 4206 3654
rect 4146 3554 4156 3594
rect 4196 3554 4206 3594
rect 3282 3454 3292 3494
rect 3332 3454 3342 3494
rect 3282 3438 3342 3454
rect 4146 3494 4206 3554
rect 4146 3454 4156 3494
rect 4196 3454 4206 3494
rect 4146 3438 4206 3454
rect 4290 3794 4350 3810
rect 4290 3754 4300 3794
rect 4340 3754 4350 3794
rect 4290 3694 4350 3754
rect 4290 3654 4300 3694
rect 4340 3654 4350 3694
rect 4290 3594 4350 3654
rect 4290 3554 4300 3594
rect 4340 3554 4350 3594
rect 4290 3494 4350 3554
rect 4290 3454 4300 3494
rect 4340 3454 4350 3494
rect 4290 3438 4350 3454
rect 4434 3794 4494 3810
rect 4434 3754 4444 3794
rect 4484 3754 4494 3794
rect 4434 3694 4494 3754
rect 4434 3654 4444 3694
rect 4484 3654 4494 3694
rect 4434 3594 4494 3654
rect 4434 3554 4444 3594
rect 4484 3554 4494 3594
rect 4434 3494 4494 3554
rect 4434 3454 4444 3494
rect 4484 3454 4494 3494
rect 4434 3438 4494 3454
rect 4722 3794 4782 3810
rect 4722 3754 4732 3794
rect 4772 3754 4782 3794
rect 4722 3694 4782 3754
rect 4722 3654 4732 3694
rect 4772 3654 4782 3694
rect 4722 3594 4782 3654
rect 4722 3554 4732 3594
rect 4772 3554 4782 3594
rect 4722 3494 4782 3554
rect 4722 3454 4732 3494
rect 4772 3454 4782 3494
rect 4722 3438 4782 3454
rect 4866 3794 4926 3810
rect 4866 3754 4876 3794
rect 4916 3754 4926 3794
rect 4866 3694 4926 3754
rect 4866 3654 4876 3694
rect 4916 3654 4926 3694
rect 4866 3594 4926 3654
rect 4866 3554 4876 3594
rect 4916 3554 4926 3594
rect 4866 3494 4926 3554
rect 4866 3454 4876 3494
rect 4916 3454 4926 3494
rect 4866 3438 4926 3454
rect 5010 3794 5070 3810
rect 5010 3754 5020 3794
rect 5060 3754 5070 3794
rect 5010 3694 5070 3754
rect 5010 3654 5020 3694
rect 5060 3654 5070 3694
rect 5010 3594 5070 3654
rect 5010 3554 5020 3594
rect 5060 3554 5070 3594
rect 5010 3494 5070 3554
rect 5010 3454 5020 3494
rect 5060 3454 5070 3494
rect 5010 3438 5070 3454
rect 5298 3794 5358 3810
rect 5298 3754 5308 3794
rect 5348 3754 5358 3794
rect 5298 3694 5358 3754
rect 5298 3654 5308 3694
rect 5348 3654 5358 3694
rect 5298 3594 5358 3654
rect 5298 3554 5308 3594
rect 5348 3554 5358 3594
rect 5298 3494 5358 3554
rect 5298 3454 5308 3494
rect 5348 3454 5358 3494
rect 5298 3438 5358 3454
rect 5442 3794 5502 3810
rect 5442 3754 5452 3794
rect 5492 3754 5502 3794
rect 5442 3694 5502 3754
rect 5442 3654 5452 3694
rect 5492 3654 5502 3694
rect 5442 3594 5502 3654
rect 5442 3554 5452 3594
rect 5492 3554 5502 3594
rect 5442 3494 5502 3554
rect 5442 3454 5452 3494
rect 5492 3454 5502 3494
rect 5442 3438 5502 3454
rect 5586 3794 5646 3810
rect 5586 3754 5596 3794
rect 5636 3754 5646 3794
rect 5586 3694 5646 3754
rect 5586 3654 5596 3694
rect 5636 3654 5646 3694
rect 5586 3594 5646 3654
rect 5586 3554 5596 3594
rect 5636 3554 5646 3594
rect 5586 3494 5646 3554
rect 5586 3454 5596 3494
rect 5636 3454 5646 3494
rect 5586 3438 5646 3454
rect 5874 3794 5934 3810
rect 5874 3754 5884 3794
rect 5924 3754 5934 3794
rect 5874 3694 5934 3754
rect 5874 3654 5884 3694
rect 5924 3654 5934 3694
rect 5874 3594 5934 3654
rect 5874 3554 5884 3594
rect 5924 3554 5934 3594
rect 5874 3494 5934 3554
rect 5874 3454 5884 3494
rect 5924 3454 5934 3494
rect 5874 3438 5934 3454
rect 6018 3794 6078 3810
rect 6018 3754 6028 3794
rect 6068 3754 6078 3794
rect 6018 3694 6078 3754
rect 6018 3654 6028 3694
rect 6068 3654 6078 3694
rect 6018 3594 6078 3654
rect 6018 3554 6028 3594
rect 6068 3554 6078 3594
rect 6018 3494 6078 3554
rect 6018 3454 6028 3494
rect 6068 3454 6078 3494
rect 6018 3438 6078 3454
rect 6162 3794 6222 3810
rect 6162 3754 6172 3794
rect 6212 3754 6222 3794
rect 6162 3694 6222 3754
rect 6162 3654 6172 3694
rect 6212 3654 6222 3694
rect 6162 3594 6222 3654
rect 6162 3554 6172 3594
rect 6212 3554 6222 3594
rect 6162 3494 6222 3554
rect 6162 3454 6172 3494
rect 6212 3454 6222 3494
rect 6162 3438 6222 3454
rect 6450 3794 6510 3810
rect 6450 3754 6460 3794
rect 6500 3754 6510 3794
rect 6450 3694 6510 3754
rect 6450 3654 6460 3694
rect 6500 3654 6510 3694
rect 6450 3594 6510 3654
rect 6450 3554 6460 3594
rect 6500 3554 6510 3594
rect 6450 3494 6510 3554
rect 6450 3454 6460 3494
rect 6500 3454 6510 3494
rect 6450 3438 6510 3454
rect 6594 3794 6654 3810
rect 6594 3754 6604 3794
rect 6644 3754 6654 3794
rect 6594 3694 6654 3754
rect 6594 3654 6604 3694
rect 6644 3654 6654 3694
rect 6594 3594 6654 3654
rect 6594 3554 6604 3594
rect 6644 3554 6654 3594
rect 6594 3494 6654 3554
rect 6594 3454 6604 3494
rect 6644 3454 6654 3494
rect 6594 3438 6654 3454
rect 6738 3794 6798 3810
rect 6738 3754 6748 3794
rect 6788 3754 6798 3794
rect 6738 3694 6798 3754
rect 7602 3794 7662 3810
rect 7602 3754 7612 3794
rect 7652 3754 7662 3794
rect 6738 3654 6748 3694
rect 6788 3654 6798 3694
rect 6738 3594 6798 3654
rect 6738 3554 6748 3594
rect 6788 3554 6798 3594
rect 6738 3494 6798 3554
rect 7026 3704 7086 3728
rect 7026 3552 7036 3704
rect 7076 3552 7086 3704
rect 7026 3528 7086 3552
rect 7170 3704 7230 3728
rect 7170 3552 7180 3704
rect 7220 3552 7230 3704
rect 7170 3528 7230 3552
rect 7314 3704 7374 3728
rect 7314 3552 7324 3704
rect 7364 3552 7374 3704
rect 7314 3528 7374 3552
rect 7602 3694 7662 3754
rect 7602 3654 7612 3694
rect 7652 3654 7662 3694
rect 7602 3594 7662 3654
rect 7602 3554 7612 3594
rect 7652 3554 7662 3594
rect 6738 3454 6748 3494
rect 6788 3454 6798 3494
rect 6738 3438 6798 3454
rect 7602 3494 7662 3554
rect 7602 3454 7612 3494
rect 7652 3454 7662 3494
rect 7602 3438 7662 3454
rect 7746 3794 7806 3810
rect 7746 3754 7756 3794
rect 7796 3754 7806 3794
rect 7746 3694 7806 3754
rect 7746 3654 7756 3694
rect 7796 3654 7806 3694
rect 7746 3594 7806 3654
rect 7746 3554 7756 3594
rect 7796 3554 7806 3594
rect 7746 3494 7806 3554
rect 7746 3454 7756 3494
rect 7796 3454 7806 3494
rect 7746 3438 7806 3454
rect 7890 3794 7950 3810
rect 7890 3754 7900 3794
rect 7940 3754 7950 3794
rect 7890 3694 7950 3754
rect 7890 3654 7900 3694
rect 7940 3654 7950 3694
rect 7890 3594 7950 3654
rect 7890 3554 7900 3594
rect 7940 3554 7950 3594
rect 7890 3494 7950 3554
rect 7890 3454 7900 3494
rect 7940 3454 7950 3494
rect 7890 3438 7950 3454
rect 8178 3794 8238 3810
rect 8178 3754 8188 3794
rect 8228 3754 8238 3794
rect 8178 3694 8238 3754
rect 8178 3654 8188 3694
rect 8228 3654 8238 3694
rect 8178 3594 8238 3654
rect 8178 3554 8188 3594
rect 8228 3554 8238 3594
rect 8178 3494 8238 3554
rect 8178 3454 8188 3494
rect 8228 3454 8238 3494
rect 8178 3438 8238 3454
rect 8322 3794 8382 3810
rect 8322 3754 8332 3794
rect 8372 3754 8382 3794
rect 8322 3694 8382 3754
rect 8322 3654 8332 3694
rect 8372 3654 8382 3694
rect 8322 3594 8382 3654
rect 8322 3554 8332 3594
rect 8372 3554 8382 3594
rect 8322 3494 8382 3554
rect 8322 3454 8332 3494
rect 8372 3454 8382 3494
rect 8322 3438 8382 3454
rect 8466 3794 8526 3810
rect 8466 3754 8476 3794
rect 8516 3754 8526 3794
rect 8466 3694 8526 3754
rect 8466 3654 8476 3694
rect 8516 3654 8526 3694
rect 8466 3594 8526 3654
rect 8466 3554 8476 3594
rect 8516 3554 8526 3594
rect 8466 3494 8526 3554
rect 8466 3454 8476 3494
rect 8516 3454 8526 3494
rect 8466 3438 8526 3454
rect 8754 3794 8814 3810
rect 8754 3754 8764 3794
rect 8804 3754 8814 3794
rect 8754 3694 8814 3754
rect 8754 3654 8764 3694
rect 8804 3654 8814 3694
rect 8754 3594 8814 3654
rect 8754 3554 8764 3594
rect 8804 3554 8814 3594
rect 8754 3494 8814 3554
rect 8754 3454 8764 3494
rect 8804 3454 8814 3494
rect 8754 3438 8814 3454
rect 8898 3794 8958 3810
rect 8898 3754 8908 3794
rect 8948 3754 8958 3794
rect 8898 3694 8958 3754
rect 8898 3654 8908 3694
rect 8948 3654 8958 3694
rect 8898 3594 8958 3654
rect 8898 3554 8908 3594
rect 8948 3554 8958 3594
rect 8898 3494 8958 3554
rect 8898 3454 8908 3494
rect 8948 3454 8958 3494
rect 8898 3438 8958 3454
rect 9042 3794 9102 3810
rect 9042 3754 9052 3794
rect 9092 3754 9102 3794
rect 9042 3694 9102 3754
rect 9042 3654 9052 3694
rect 9092 3654 9102 3694
rect 9042 3594 9102 3654
rect 9042 3554 9052 3594
rect 9092 3554 9102 3594
rect 9042 3494 9102 3554
rect 9042 3454 9052 3494
rect 9092 3454 9102 3494
rect 9042 3438 9102 3454
rect 9330 3794 9390 3810
rect 9330 3754 9340 3794
rect 9380 3754 9390 3794
rect 9330 3694 9390 3754
rect 9330 3654 9340 3694
rect 9380 3654 9390 3694
rect 9330 3594 9390 3654
rect 9330 3554 9340 3594
rect 9380 3554 9390 3594
rect 9330 3494 9390 3554
rect 9330 3454 9340 3494
rect 9380 3454 9390 3494
rect 9330 3438 9390 3454
rect 9474 3794 9534 3810
rect 9474 3754 9484 3794
rect 9524 3754 9534 3794
rect 9474 3694 9534 3754
rect 9474 3654 9484 3694
rect 9524 3654 9534 3694
rect 9474 3594 9534 3654
rect 9474 3554 9484 3594
rect 9524 3554 9534 3594
rect 9474 3494 9534 3554
rect 9474 3454 9484 3494
rect 9524 3454 9534 3494
rect 9474 3438 9534 3454
rect 9618 3794 9678 3810
rect 9618 3754 9628 3794
rect 9668 3754 9678 3794
rect 9618 3694 9678 3754
rect 9618 3654 9628 3694
rect 9668 3654 9678 3694
rect 9618 3594 9678 3654
rect 9618 3554 9628 3594
rect 9668 3554 9678 3594
rect 9618 3494 9678 3554
rect 9618 3454 9628 3494
rect 9668 3454 9678 3494
rect 9618 3438 9678 3454
rect 10194 3794 10254 3810
rect 10194 3754 10204 3794
rect 10244 3754 10254 3794
rect 10194 3694 10254 3754
rect 10194 3654 10204 3694
rect 10244 3654 10254 3694
rect 10194 3594 10254 3654
rect 10194 3554 10204 3594
rect 10244 3554 10254 3594
rect 10194 3494 10254 3554
rect 10194 3454 10204 3494
rect 10244 3454 10254 3494
rect 10194 3438 10254 3454
rect 10338 3794 10398 3810
rect 10338 3754 10348 3794
rect 10388 3754 10398 3794
rect 10338 3694 10398 3754
rect 10338 3654 10348 3694
rect 10388 3654 10398 3694
rect 10338 3594 10398 3654
rect 10338 3554 10348 3594
rect 10388 3554 10398 3594
rect 10338 3494 10398 3554
rect 10338 3454 10348 3494
rect 10388 3454 10398 3494
rect 10338 3438 10398 3454
rect 10482 3794 10542 3810
rect 10482 3754 10492 3794
rect 10532 3754 10542 3794
rect 10482 3694 10542 3754
rect 10482 3654 10492 3694
rect 10532 3654 10542 3694
rect 10482 3594 10542 3654
rect 10482 3554 10492 3594
rect 10532 3554 10542 3594
rect 10482 3494 10542 3554
rect 10482 3454 10492 3494
rect 10532 3454 10542 3494
rect 10482 3438 10542 3454
rect 10770 3794 10830 3810
rect 10770 3754 10780 3794
rect 10820 3754 10830 3794
rect 10770 3694 10830 3754
rect 10770 3654 10780 3694
rect 10820 3654 10830 3694
rect 10770 3594 10830 3654
rect 10770 3554 10780 3594
rect 10820 3554 10830 3594
rect 10770 3494 10830 3554
rect 10770 3454 10780 3494
rect 10820 3454 10830 3494
rect 10770 3438 10830 3454
rect 10914 3794 10974 3810
rect 10914 3754 10924 3794
rect 10964 3754 10974 3794
rect 10914 3694 10974 3754
rect 10914 3654 10924 3694
rect 10964 3654 10974 3694
rect 10914 3594 10974 3654
rect 10914 3554 10924 3594
rect 10964 3554 10974 3594
rect 10914 3494 10974 3554
rect 10914 3454 10924 3494
rect 10964 3454 10974 3494
rect 10914 3438 10974 3454
rect 11058 3794 11118 3810
rect 11058 3754 11068 3794
rect 11108 3754 11118 3794
rect 11058 3694 11118 3754
rect 11922 3794 11982 3810
rect 11922 3754 11932 3794
rect 11972 3754 11982 3794
rect 11058 3654 11068 3694
rect 11108 3654 11118 3694
rect 11058 3594 11118 3654
rect 11058 3554 11068 3594
rect 11108 3554 11118 3594
rect 11058 3494 11118 3554
rect 11346 3704 11406 3728
rect 11346 3552 11356 3704
rect 11396 3552 11406 3704
rect 11346 3528 11406 3552
rect 11490 3704 11550 3728
rect 11490 3552 11500 3704
rect 11540 3552 11550 3704
rect 11490 3528 11550 3552
rect 11634 3704 11694 3728
rect 11634 3552 11644 3704
rect 11684 3552 11694 3704
rect 11634 3528 11694 3552
rect 11922 3694 11982 3754
rect 11922 3654 11932 3694
rect 11972 3654 11982 3694
rect 11922 3594 11982 3654
rect 11922 3554 11932 3594
rect 11972 3554 11982 3594
rect 11058 3454 11068 3494
rect 11108 3454 11118 3494
rect 11058 3438 11118 3454
rect 11922 3494 11982 3554
rect 11922 3454 11932 3494
rect 11972 3454 11982 3494
rect 11922 3438 11982 3454
rect 12066 3794 12126 3810
rect 12066 3754 12076 3794
rect 12116 3754 12126 3794
rect 12066 3694 12126 3754
rect 12066 3654 12076 3694
rect 12116 3654 12126 3694
rect 12066 3594 12126 3654
rect 12066 3554 12076 3594
rect 12116 3554 12126 3594
rect 12066 3494 12126 3554
rect 12066 3454 12076 3494
rect 12116 3454 12126 3494
rect 12066 3438 12126 3454
rect 12210 3794 12270 3810
rect 12210 3754 12220 3794
rect 12260 3754 12270 3794
rect 12210 3694 12270 3754
rect 12210 3654 12220 3694
rect 12260 3654 12270 3694
rect 12210 3594 12270 3654
rect 12210 3554 12220 3594
rect 12260 3554 12270 3594
rect 12210 3494 12270 3554
rect 12210 3454 12220 3494
rect 12260 3454 12270 3494
rect 12210 3438 12270 3454
rect 12498 3794 12558 3810
rect 12498 3754 12508 3794
rect 12548 3754 12558 3794
rect 12498 3694 12558 3754
rect 12498 3654 12508 3694
rect 12548 3654 12558 3694
rect 12498 3594 12558 3654
rect 12498 3554 12508 3594
rect 12548 3554 12558 3594
rect 12498 3494 12558 3554
rect 12498 3454 12508 3494
rect 12548 3454 12558 3494
rect 12498 3438 12558 3454
rect 12642 3794 12702 3810
rect 12642 3754 12652 3794
rect 12692 3754 12702 3794
rect 12642 3694 12702 3754
rect 12642 3654 12652 3694
rect 12692 3654 12702 3694
rect 12642 3594 12702 3654
rect 12642 3554 12652 3594
rect 12692 3554 12702 3594
rect 12642 3494 12702 3554
rect 12642 3454 12652 3494
rect 12692 3454 12702 3494
rect 12642 3438 12702 3454
rect 12786 3794 12846 3810
rect 12786 3754 12796 3794
rect 12836 3754 12846 3794
rect 12786 3694 12846 3754
rect 12786 3654 12796 3694
rect 12836 3654 12846 3694
rect 12786 3594 12846 3654
rect 12786 3554 12796 3594
rect 12836 3554 12846 3594
rect 12786 3494 12846 3554
rect 12786 3454 12796 3494
rect 12836 3454 12846 3494
rect 12786 3438 12846 3454
rect 13650 3794 13710 3810
rect 13650 3754 13660 3794
rect 13700 3754 13710 3794
rect 13650 3694 13710 3754
rect 13650 3654 13660 3694
rect 13700 3654 13710 3694
rect 13650 3594 13710 3654
rect 13650 3554 13660 3594
rect 13700 3554 13710 3594
rect 13650 3494 13710 3554
rect 13650 3454 13660 3494
rect 13700 3454 13710 3494
rect 13650 3438 13710 3454
rect 13794 3794 13854 3810
rect 13794 3754 13804 3794
rect 13844 3754 13854 3794
rect 13794 3694 13854 3754
rect 13794 3654 13804 3694
rect 13844 3654 13854 3694
rect 13794 3594 13854 3654
rect 13794 3554 13804 3594
rect 13844 3554 13854 3594
rect 13794 3494 13854 3554
rect 13794 3454 13804 3494
rect 13844 3454 13854 3494
rect 13794 3438 13854 3454
rect 13938 3794 13998 3810
rect 13938 3754 13948 3794
rect 13988 3754 13998 3794
rect 13938 3694 13998 3754
rect 13938 3654 13948 3694
rect 13988 3654 13998 3694
rect 13938 3594 13998 3654
rect 13938 3554 13948 3594
rect 13988 3554 13998 3594
rect 13938 3494 13998 3554
rect 13938 3454 13948 3494
rect 13988 3454 13998 3494
rect 13938 3438 13998 3454
rect 14226 3794 14286 3810
rect 14226 3754 14236 3794
rect 14276 3754 14286 3794
rect 14226 3694 14286 3754
rect 14226 3654 14236 3694
rect 14276 3654 14286 3694
rect 14226 3594 14286 3654
rect 14226 3554 14236 3594
rect 14276 3554 14286 3594
rect 14226 3494 14286 3554
rect 14226 3454 14236 3494
rect 14276 3454 14286 3494
rect 14226 3438 14286 3454
rect 14370 3794 14430 3810
rect 14370 3754 14380 3794
rect 14420 3754 14430 3794
rect 14370 3694 14430 3754
rect 14370 3654 14380 3694
rect 14420 3654 14430 3694
rect 14370 3594 14430 3654
rect 14370 3554 14380 3594
rect 14420 3554 14430 3594
rect 14370 3494 14430 3554
rect 14370 3454 14380 3494
rect 14420 3454 14430 3494
rect 14370 3438 14430 3454
rect 14514 3794 14574 3810
rect 14514 3754 14524 3794
rect 14564 3754 14574 3794
rect 14514 3694 14574 3754
rect 14514 3654 14524 3694
rect 14564 3654 14574 3694
rect 14514 3594 14574 3654
rect 14514 3554 14524 3594
rect 14564 3554 14574 3594
rect 14514 3494 14574 3554
rect 14514 3454 14524 3494
rect 14564 3454 14574 3494
rect 14514 3438 14574 3454
rect 14802 3794 14862 3810
rect 14802 3754 14812 3794
rect 14852 3754 14862 3794
rect 14802 3694 14862 3754
rect 14802 3654 14812 3694
rect 14852 3654 14862 3694
rect 14802 3594 14862 3654
rect 14802 3554 14812 3594
rect 14852 3554 14862 3594
rect 14802 3494 14862 3554
rect 14802 3454 14812 3494
rect 14852 3454 14862 3494
rect 14802 3438 14862 3454
rect 14946 3794 15006 3810
rect 14946 3754 14956 3794
rect 14996 3754 15006 3794
rect 14946 3694 15006 3754
rect 14946 3654 14956 3694
rect 14996 3654 15006 3694
rect 14946 3594 15006 3654
rect 14946 3554 14956 3594
rect 14996 3554 15006 3594
rect 14946 3494 15006 3554
rect 14946 3454 14956 3494
rect 14996 3454 15006 3494
rect 14946 3438 15006 3454
rect 15090 3794 15150 3810
rect 15090 3754 15100 3794
rect 15140 3754 15150 3794
rect 15090 3694 15150 3754
rect 16530 3794 16590 3810
rect 16530 3754 16540 3794
rect 16580 3754 16590 3794
rect 15090 3654 15100 3694
rect 15140 3654 15150 3694
rect 15090 3594 15150 3654
rect 15090 3554 15100 3594
rect 15140 3554 15150 3594
rect 15090 3494 15150 3554
rect 15378 3704 15438 3728
rect 15378 3552 15388 3704
rect 15428 3552 15438 3704
rect 15378 3528 15438 3552
rect 15522 3704 15582 3728
rect 15522 3552 15532 3704
rect 15572 3552 15582 3704
rect 15522 3528 15582 3552
rect 15666 3704 15726 3728
rect 15666 3552 15676 3704
rect 15716 3552 15726 3704
rect 15666 3528 15726 3552
rect 15954 3704 16014 3728
rect 15954 3552 15964 3704
rect 16004 3552 16014 3704
rect 15954 3528 16014 3552
rect 16098 3704 16158 3728
rect 16098 3552 16108 3704
rect 16148 3552 16158 3704
rect 16098 3528 16158 3552
rect 16242 3704 16302 3728
rect 16242 3552 16252 3704
rect 16292 3552 16302 3704
rect 16242 3528 16302 3552
rect 16530 3694 16590 3754
rect 16530 3654 16540 3694
rect 16580 3654 16590 3694
rect 16530 3594 16590 3654
rect 16530 3554 16540 3594
rect 16580 3554 16590 3594
rect 15090 3454 15100 3494
rect 15140 3454 15150 3494
rect 15090 3438 15150 3454
rect 16530 3494 16590 3554
rect 16530 3454 16540 3494
rect 16580 3454 16590 3494
rect 16530 3438 16590 3454
rect 16674 3794 16734 3810
rect 16674 3754 16684 3794
rect 16724 3754 16734 3794
rect 16674 3694 16734 3754
rect 16674 3654 16684 3694
rect 16724 3654 16734 3694
rect 16674 3594 16734 3654
rect 16674 3554 16684 3594
rect 16724 3554 16734 3594
rect 16674 3494 16734 3554
rect 16674 3454 16684 3494
rect 16724 3454 16734 3494
rect 16674 3438 16734 3454
rect 16818 3794 16878 3810
rect 16818 3754 16828 3794
rect 16868 3754 16878 3794
rect 16818 3694 16878 3754
rect 16818 3654 16828 3694
rect 16868 3654 16878 3694
rect 16818 3594 16878 3654
rect 16818 3554 16828 3594
rect 16868 3554 16878 3594
rect 16818 3494 16878 3554
rect 16818 3454 16828 3494
rect 16868 3454 16878 3494
rect 16818 3438 16878 3454
rect 16962 3794 17022 3810
rect 16962 3754 16972 3794
rect 17012 3754 17022 3794
rect 16962 3694 17022 3754
rect 16962 3654 16972 3694
rect 17012 3654 17022 3694
rect 16962 3594 17022 3654
rect 16962 3554 16972 3594
rect 17012 3554 17022 3594
rect 16962 3494 17022 3554
rect 16962 3454 16972 3494
rect 17012 3454 17022 3494
rect 16962 3438 17022 3454
rect 17106 3794 17166 3810
rect 17106 3754 17116 3794
rect 17156 3754 17166 3794
rect 17106 3694 17166 3754
rect 17106 3654 17116 3694
rect 17156 3654 17166 3694
rect 17106 3594 17166 3654
rect 17106 3554 17116 3594
rect 17156 3554 17166 3594
rect 17106 3494 17166 3554
rect 17106 3454 17116 3494
rect 17156 3454 17166 3494
rect 17106 3438 17166 3454
rect 17250 3794 17310 3810
rect 17250 3754 17260 3794
rect 17300 3754 17310 3794
rect 17250 3694 17310 3754
rect 17250 3654 17260 3694
rect 17300 3654 17310 3694
rect 17250 3594 17310 3654
rect 17250 3554 17260 3594
rect 17300 3554 17310 3594
rect 17250 3494 17310 3554
rect 17250 3454 17260 3494
rect 17300 3454 17310 3494
rect 17250 3438 17310 3454
rect 17394 3794 17454 3810
rect 17394 3754 17404 3794
rect 17444 3754 17454 3794
rect 17394 3694 17454 3754
rect 17394 3654 17404 3694
rect 17444 3654 17454 3694
rect 17394 3594 17454 3654
rect 17394 3554 17404 3594
rect 17444 3554 17454 3594
rect 17394 3494 17454 3554
rect 17394 3454 17404 3494
rect 17444 3454 17454 3494
rect 17394 3438 17454 3454
rect 17538 3794 17598 3810
rect 17538 3754 17548 3794
rect 17588 3754 17598 3794
rect 17538 3694 17598 3754
rect 17538 3654 17548 3694
rect 17588 3654 17598 3694
rect 17538 3594 17598 3654
rect 17538 3554 17548 3594
rect 17588 3554 17598 3594
rect 17538 3494 17598 3554
rect 17538 3454 17548 3494
rect 17588 3454 17598 3494
rect 17538 3438 17598 3454
rect 17682 3794 17742 3810
rect 17682 3754 17692 3794
rect 17732 3754 17742 3794
rect 17682 3694 17742 3754
rect 17682 3654 17692 3694
rect 17732 3654 17742 3694
rect 17682 3594 17742 3654
rect 17682 3554 17692 3594
rect 17732 3554 17742 3594
rect 17682 3494 17742 3554
rect 17682 3454 17692 3494
rect 17732 3454 17742 3494
rect 17682 3438 17742 3454
rect 17826 3794 17886 3810
rect 17826 3754 17836 3794
rect 17876 3754 17886 3794
rect 17826 3694 17886 3754
rect 17826 3654 17836 3694
rect 17876 3654 17886 3694
rect 17826 3594 17886 3654
rect 17826 3554 17836 3594
rect 17876 3554 17886 3594
rect 17826 3494 17886 3554
rect 17826 3454 17836 3494
rect 17876 3454 17886 3494
rect 17826 3438 17886 3454
rect 17970 3794 18030 3810
rect 17970 3754 17980 3794
rect 18020 3754 18030 3794
rect 17970 3694 18030 3754
rect 17970 3654 17980 3694
rect 18020 3654 18030 3694
rect 17970 3594 18030 3654
rect 17970 3554 17980 3594
rect 18020 3554 18030 3594
rect 17970 3494 18030 3554
rect 17970 3454 17980 3494
rect 18020 3454 18030 3494
rect 17970 3438 18030 3454
rect 18114 3794 18174 3810
rect 18114 3754 18124 3794
rect 18164 3754 18174 3794
rect 18114 3694 18174 3754
rect 18114 3654 18124 3694
rect 18164 3654 18174 3694
rect 18114 3594 18174 3654
rect 18114 3554 18124 3594
rect 18164 3554 18174 3594
rect 18114 3494 18174 3554
rect 18114 3454 18124 3494
rect 18164 3454 18174 3494
rect 18114 3438 18174 3454
rect 18258 3794 18318 3810
rect 18258 3754 18268 3794
rect 18308 3754 18318 3794
rect 18258 3694 18318 3754
rect 18258 3654 18268 3694
rect 18308 3654 18318 3694
rect 18258 3594 18318 3654
rect 18258 3554 18268 3594
rect 18308 3554 18318 3594
rect 18258 3494 18318 3554
rect 18258 3454 18268 3494
rect 18308 3454 18318 3494
rect 18258 3438 18318 3454
rect 18402 3794 18462 3810
rect 18402 3754 18412 3794
rect 18452 3754 18462 3794
rect 18402 3694 18462 3754
rect 18402 3654 18412 3694
rect 18452 3654 18462 3694
rect 18402 3594 18462 3654
rect 18402 3554 18412 3594
rect 18452 3554 18462 3594
rect 18402 3494 18462 3554
rect 18402 3454 18412 3494
rect 18452 3454 18462 3494
rect 18402 3438 18462 3454
rect 18546 3794 18606 3810
rect 18546 3754 18556 3794
rect 18596 3754 18606 3794
rect 18546 3694 18606 3754
rect 18546 3654 18556 3694
rect 18596 3654 18606 3694
rect 18546 3594 18606 3654
rect 18546 3554 18556 3594
rect 18596 3554 18606 3594
rect 18546 3494 18606 3554
rect 18546 3454 18556 3494
rect 18596 3454 18606 3494
rect 18546 3438 18606 3454
rect 18690 3794 18750 3810
rect 18690 3754 18700 3794
rect 18740 3754 18750 3794
rect 18690 3694 18750 3754
rect 18690 3654 18700 3694
rect 18740 3654 18750 3694
rect 18690 3594 18750 3654
rect 18690 3554 18700 3594
rect 18740 3554 18750 3594
rect 18690 3494 18750 3554
rect 18690 3454 18700 3494
rect 18740 3454 18750 3494
rect 18690 3438 18750 3454
rect 18834 3794 18894 3810
rect 18834 3754 18844 3794
rect 18884 3754 18894 3794
rect 18834 3694 18894 3754
rect 18834 3654 18844 3694
rect 18884 3654 18894 3694
rect 18834 3594 18894 3654
rect 18834 3554 18844 3594
rect 18884 3554 18894 3594
rect 18834 3494 18894 3554
rect 18834 3454 18844 3494
rect 18884 3454 18894 3494
rect 18834 3438 18894 3454
rect 18978 3794 19038 3810
rect 18978 3754 18988 3794
rect 19028 3754 19038 3794
rect 18978 3694 19038 3754
rect 18978 3654 18988 3694
rect 19028 3654 19038 3694
rect 18978 3594 19038 3654
rect 18978 3554 18988 3594
rect 19028 3554 19038 3594
rect 18978 3494 19038 3554
rect 18978 3454 18988 3494
rect 19028 3454 19038 3494
rect 18978 3438 19038 3454
rect 19122 3794 19182 3810
rect 19122 3754 19132 3794
rect 19172 3754 19182 3794
rect 19122 3694 19182 3754
rect 19122 3654 19132 3694
rect 19172 3654 19182 3694
rect 19122 3594 19182 3654
rect 19122 3554 19132 3594
rect 19172 3554 19182 3594
rect 19122 3494 19182 3554
rect 19122 3454 19132 3494
rect 19172 3454 19182 3494
rect 19122 3438 19182 3454
rect 19266 3794 19326 3810
rect 19266 3754 19276 3794
rect 19316 3754 19326 3794
rect 19266 3694 19326 3754
rect 19266 3654 19276 3694
rect 19316 3654 19326 3694
rect 19266 3594 19326 3654
rect 19266 3554 19276 3594
rect 19316 3554 19326 3594
rect 19266 3494 19326 3554
rect 19266 3454 19276 3494
rect 19316 3454 19326 3494
rect 19266 3438 19326 3454
rect 19410 3794 19470 3810
rect 19410 3754 19420 3794
rect 19460 3754 19470 3794
rect 19410 3694 19470 3754
rect 19410 3654 19420 3694
rect 19460 3654 19470 3694
rect 19410 3594 19470 3654
rect 19410 3554 19420 3594
rect 19460 3554 19470 3594
rect 19410 3494 19470 3554
rect 19410 3454 19420 3494
rect 19460 3454 19470 3494
rect 19410 3438 19470 3454
rect 19554 3794 19614 3810
rect 19554 3754 19564 3794
rect 19604 3754 19614 3794
rect 19554 3694 19614 3754
rect 19554 3654 19564 3694
rect 19604 3654 19614 3694
rect 19554 3594 19614 3654
rect 19554 3554 19564 3594
rect 19604 3554 19614 3594
rect 19554 3494 19614 3554
rect 19554 3454 19564 3494
rect 19604 3454 19614 3494
rect 19554 3438 19614 3454
rect 19698 3794 19758 3810
rect 19698 3754 19708 3794
rect 19748 3754 19758 3794
rect 19698 3694 19758 3754
rect 19698 3654 19708 3694
rect 19748 3654 19758 3694
rect 19698 3594 19758 3654
rect 19698 3554 19708 3594
rect 19748 3554 19758 3594
rect 19698 3494 19758 3554
rect 19698 3454 19708 3494
rect 19748 3454 19758 3494
rect 19698 3438 19758 3454
rect 19842 3794 19902 3810
rect 19842 3754 19852 3794
rect 19892 3754 19902 3794
rect 19842 3694 19902 3754
rect 19842 3654 19852 3694
rect 19892 3654 19902 3694
rect 19842 3594 19902 3654
rect 19842 3554 19852 3594
rect 19892 3554 19902 3594
rect 19842 3494 19902 3554
rect 19842 3454 19852 3494
rect 19892 3454 19902 3494
rect 19842 3438 19902 3454
rect 19986 3794 20046 3810
rect 19986 3754 19996 3794
rect 20036 3754 20046 3794
rect 19986 3694 20046 3754
rect 19986 3654 19996 3694
rect 20036 3654 20046 3694
rect 19986 3594 20046 3654
rect 19986 3554 19996 3594
rect 20036 3554 20046 3594
rect 19986 3494 20046 3554
rect 19986 3454 19996 3494
rect 20036 3454 20046 3494
rect 19986 3438 20046 3454
rect 778 3329 952 3348
rect 778 3295 790 3329
rect 824 3295 898 3329
rect 932 3295 952 3329
rect 778 3276 952 3295
rect 1354 3329 1528 3348
rect 1354 3295 1366 3329
rect 1400 3295 1474 3329
rect 1508 3295 1528 3329
rect 1354 3276 1528 3295
rect 1930 3329 2104 3348
rect 1930 3295 1942 3329
rect 1976 3295 2050 3329
rect 2084 3295 2104 3329
rect 1930 3276 2104 3295
rect 2506 3329 2680 3348
rect 2506 3295 2518 3329
rect 2552 3295 2626 3329
rect 2660 3295 2680 3329
rect 2506 3276 2680 3295
rect 3080 3329 3254 3348
rect 3080 3295 3100 3329
rect 3134 3295 3208 3329
rect 3242 3295 3254 3329
rect 3080 3276 3254 3295
rect 4232 3329 4406 3348
rect 4232 3295 4252 3329
rect 4286 3295 4360 3329
rect 4394 3295 4406 3329
rect 4232 3276 4406 3295
rect 4808 3329 4982 3348
rect 4808 3295 4828 3329
rect 4862 3295 4936 3329
rect 4970 3295 4982 3329
rect 4808 3276 4982 3295
rect 5384 3329 5558 3348
rect 5384 3295 5404 3329
rect 5438 3295 5512 3329
rect 5546 3295 5558 3329
rect 5384 3276 5558 3295
rect 5960 3329 6134 3348
rect 5960 3295 5980 3329
rect 6014 3295 6088 3329
rect 6122 3295 6134 3329
rect 5960 3276 6134 3295
rect 6446 3330 6536 3348
rect 6446 3294 6468 3330
rect 6504 3294 6536 3330
rect 6446 3276 6536 3294
rect 6710 3330 6800 3348
rect 6710 3294 6752 3330
rect 6788 3294 6800 3330
rect 6710 3276 6800 3294
rect 7688 3329 7862 3348
rect 7688 3295 7708 3329
rect 7742 3295 7816 3329
rect 7850 3295 7862 3329
rect 7688 3276 7862 3295
rect 8264 3329 8438 3348
rect 8264 3295 8284 3329
rect 8318 3295 8392 3329
rect 8426 3295 8438 3329
rect 8264 3276 8438 3295
rect 8840 3329 9014 3348
rect 8840 3295 8860 3329
rect 8894 3295 8968 3329
rect 9002 3295 9014 3329
rect 8840 3276 9014 3295
rect 9326 3330 9416 3348
rect 9326 3294 9348 3330
rect 9384 3294 9416 3330
rect 9326 3276 9416 3294
rect 9590 3330 9680 3348
rect 9590 3294 9632 3330
rect 9668 3294 9680 3330
rect 9590 3276 9680 3294
rect 10280 3329 10454 3348
rect 10280 3295 10300 3329
rect 10334 3295 10408 3329
rect 10442 3295 10454 3329
rect 10280 3276 10454 3295
rect 10856 3329 11030 3348
rect 10856 3295 10876 3329
rect 10910 3295 10984 3329
rect 11018 3295 11030 3329
rect 10856 3276 11030 3295
rect 12008 3329 12182 3348
rect 12008 3295 12028 3329
rect 12062 3295 12136 3329
rect 12170 3295 12182 3329
rect 12008 3276 12182 3295
rect 12584 3329 12758 3348
rect 12584 3295 12604 3329
rect 12638 3295 12712 3329
rect 12746 3295 12758 3329
rect 12584 3276 12758 3295
rect 13736 3329 13910 3348
rect 13736 3295 13756 3329
rect 13790 3295 13864 3329
rect 13898 3295 13910 3329
rect 13736 3276 13910 3295
rect 14312 3329 14486 3348
rect 14312 3295 14332 3329
rect 14366 3295 14440 3329
rect 14474 3295 14486 3329
rect 14312 3276 14486 3295
rect 14888 3329 15062 3348
rect 14888 3295 14908 3329
rect 14942 3295 15016 3329
rect 15050 3295 15062 3329
rect 14888 3276 15062 3295
rect 16618 3329 16792 3348
rect 16618 3295 16630 3329
rect 16664 3295 16738 3329
rect 16772 3295 16792 3329
rect 16618 3276 16792 3295
rect 16906 3329 17080 3348
rect 16906 3295 16918 3329
rect 16952 3295 17026 3329
rect 17060 3295 17080 3329
rect 16906 3276 17080 3295
rect 17194 3329 17368 3348
rect 17194 3295 17206 3329
rect 17240 3295 17314 3329
rect 17348 3295 17368 3329
rect 17194 3276 17368 3295
rect 17482 3329 17656 3348
rect 17482 3295 17494 3329
rect 17528 3295 17602 3329
rect 17636 3295 17656 3329
rect 17482 3276 17656 3295
rect 17770 3329 17944 3348
rect 17770 3295 17782 3329
rect 17816 3295 17890 3329
rect 17924 3295 17944 3329
rect 17770 3276 17944 3295
rect 18058 3329 18232 3348
rect 18058 3295 18070 3329
rect 18104 3295 18178 3329
rect 18212 3295 18232 3329
rect 18058 3276 18232 3295
rect 18346 3329 18520 3348
rect 18346 3295 18358 3329
rect 18392 3295 18466 3329
rect 18500 3295 18520 3329
rect 18346 3276 18520 3295
rect 18634 3329 18808 3348
rect 18634 3295 18646 3329
rect 18680 3295 18754 3329
rect 18788 3295 18808 3329
rect 18634 3276 18808 3295
rect 18922 3329 19096 3348
rect 18922 3295 18934 3329
rect 18968 3295 19042 3329
rect 19076 3295 19096 3329
rect 18922 3276 19096 3295
rect 19210 3329 19384 3348
rect 19210 3295 19222 3329
rect 19256 3295 19330 3329
rect 19364 3295 19384 3329
rect 19210 3276 19384 3295
rect 19498 3329 19672 3348
rect 19498 3295 19510 3329
rect 19544 3295 19618 3329
rect 19652 3295 19672 3329
rect 19498 3276 19672 3295
rect 19786 3329 19960 3348
rect 19786 3295 19798 3329
rect 19832 3295 19906 3329
rect 19940 3295 19960 3329
rect 19786 3276 19960 3295
rect 778 2753 952 2772
rect 778 2719 790 2753
rect 824 2719 898 2753
rect 932 2719 952 2753
rect 778 2700 952 2719
rect 1354 2753 1528 2772
rect 1354 2719 1366 2753
rect 1400 2719 1474 2753
rect 1508 2719 1528 2753
rect 1354 2700 1528 2719
rect 1930 2753 2104 2772
rect 1930 2719 1942 2753
rect 1976 2719 2050 2753
rect 2084 2719 2104 2753
rect 1930 2700 2104 2719
rect 2506 2753 2680 2772
rect 2506 2719 2518 2753
rect 2552 2719 2626 2753
rect 2660 2719 2680 2753
rect 2506 2700 2680 2719
rect 3080 2753 3254 2772
rect 3080 2719 3100 2753
rect 3134 2719 3208 2753
rect 3242 2719 3254 2753
rect 3080 2700 3254 2719
rect 4232 2753 4406 2772
rect 4232 2719 4252 2753
rect 4286 2719 4360 2753
rect 4394 2719 4406 2753
rect 4232 2700 4406 2719
rect 4808 2753 4982 2772
rect 4808 2719 4828 2753
rect 4862 2719 4936 2753
rect 4970 2719 4982 2753
rect 4808 2700 4982 2719
rect 5384 2753 5558 2772
rect 5384 2719 5404 2753
rect 5438 2719 5512 2753
rect 5546 2719 5558 2753
rect 5384 2700 5558 2719
rect 5960 2753 6134 2772
rect 5960 2719 5980 2753
rect 6014 2719 6088 2753
rect 6122 2719 6134 2753
rect 5960 2700 6134 2719
rect 6446 2754 6536 2772
rect 6446 2718 6468 2754
rect 6504 2718 6536 2754
rect 6446 2700 6536 2718
rect 6710 2754 6800 2772
rect 6710 2718 6746 2754
rect 6782 2718 6800 2754
rect 6710 2700 6800 2718
rect 7688 2753 7862 2772
rect 7688 2719 7708 2753
rect 7742 2719 7816 2753
rect 7850 2719 7862 2753
rect 7688 2700 7862 2719
rect 8264 2753 8438 2772
rect 8264 2719 8284 2753
rect 8318 2719 8392 2753
rect 8426 2719 8438 2753
rect 8264 2700 8438 2719
rect 8840 2753 9014 2772
rect 8840 2719 8860 2753
rect 8894 2719 8968 2753
rect 9002 2719 9014 2753
rect 8840 2700 9014 2719
rect 9326 2754 9416 2772
rect 9326 2718 9348 2754
rect 9384 2718 9416 2754
rect 9326 2700 9416 2718
rect 9590 2754 9680 2772
rect 9590 2718 9626 2754
rect 9662 2718 9680 2754
rect 9590 2700 9680 2718
rect 10280 2753 10454 2772
rect 10280 2719 10300 2753
rect 10334 2719 10408 2753
rect 10442 2719 10454 2753
rect 10280 2700 10454 2719
rect 10856 2753 11030 2772
rect 10856 2719 10876 2753
rect 10910 2719 10984 2753
rect 11018 2719 11030 2753
rect 10856 2700 11030 2719
rect 12008 2753 12182 2772
rect 12008 2719 12028 2753
rect 12062 2719 12136 2753
rect 12170 2719 12182 2753
rect 12008 2700 12182 2719
rect 12584 2753 12758 2772
rect 12584 2719 12604 2753
rect 12638 2719 12712 2753
rect 12746 2719 12758 2753
rect 12584 2700 12758 2719
rect 13736 2753 13910 2772
rect 13736 2719 13756 2753
rect 13790 2719 13864 2753
rect 13898 2719 13910 2753
rect 13736 2700 13910 2719
rect 14312 2753 14486 2772
rect 14312 2719 14332 2753
rect 14366 2719 14440 2753
rect 14474 2719 14486 2753
rect 14312 2700 14486 2719
rect 14888 2753 15062 2772
rect 14888 2719 14908 2753
rect 14942 2719 15016 2753
rect 15050 2719 15062 2753
rect 14888 2700 15062 2719
rect 16618 2753 16792 2772
rect 16618 2719 16630 2753
rect 16664 2719 16738 2753
rect 16772 2719 16792 2753
rect 16618 2700 16792 2719
rect 16906 2753 17080 2772
rect 16906 2719 16918 2753
rect 16952 2719 17026 2753
rect 17060 2719 17080 2753
rect 16906 2700 17080 2719
rect 17194 2753 17368 2772
rect 17194 2719 17206 2753
rect 17240 2719 17314 2753
rect 17348 2719 17368 2753
rect 17194 2700 17368 2719
rect 17482 2753 17656 2772
rect 17482 2719 17494 2753
rect 17528 2719 17602 2753
rect 17636 2719 17656 2753
rect 17482 2700 17656 2719
rect 17770 2753 17944 2772
rect 17770 2719 17782 2753
rect 17816 2719 17890 2753
rect 17924 2719 17944 2753
rect 17770 2700 17944 2719
rect 18058 2753 18232 2772
rect 18058 2719 18070 2753
rect 18104 2719 18178 2753
rect 18212 2719 18232 2753
rect 18058 2700 18232 2719
rect 18346 2753 18520 2772
rect 18346 2719 18358 2753
rect 18392 2719 18466 2753
rect 18500 2719 18520 2753
rect 18346 2700 18520 2719
rect 18634 2753 18808 2772
rect 18634 2719 18646 2753
rect 18680 2719 18754 2753
rect 18788 2719 18808 2753
rect 18634 2700 18808 2719
rect 18922 2753 19096 2772
rect 18922 2719 18934 2753
rect 18968 2719 19042 2753
rect 19076 2719 19096 2753
rect 18922 2700 19096 2719
rect 19210 2753 19384 2772
rect 19210 2719 19222 2753
rect 19256 2719 19330 2753
rect 19364 2719 19384 2753
rect 19210 2700 19384 2719
rect 19498 2753 19672 2772
rect 19498 2719 19510 2753
rect 19544 2719 19618 2753
rect 19652 2719 19672 2753
rect 19498 2700 19672 2719
rect 19786 2753 19960 2772
rect 19786 2719 19798 2753
rect 19832 2719 19906 2753
rect 19940 2719 19960 2753
rect 19786 2700 19960 2719
rect 114 2588 174 2630
rect 114 2500 124 2588
rect 164 2500 174 2588
rect 114 2458 174 2500
rect 258 2588 318 2630
rect 258 2500 268 2588
rect 308 2500 318 2588
rect 258 2458 318 2500
rect 402 2588 462 2630
rect 402 2500 412 2588
rect 452 2500 462 2588
rect 402 2458 462 2500
rect 690 2614 750 2630
rect 690 2574 700 2614
rect 740 2574 750 2614
rect 690 2514 750 2574
rect 690 2474 700 2514
rect 740 2474 750 2514
rect 690 2458 750 2474
rect 834 2614 894 2630
rect 834 2574 844 2614
rect 884 2574 894 2614
rect 834 2514 894 2574
rect 834 2474 844 2514
rect 884 2474 894 2514
rect 834 2458 894 2474
rect 978 2614 1038 2630
rect 978 2574 988 2614
rect 1028 2574 1038 2614
rect 978 2514 1038 2574
rect 978 2474 988 2514
rect 1028 2474 1038 2514
rect 978 2458 1038 2474
rect 1266 2614 1326 2630
rect 1266 2574 1276 2614
rect 1316 2574 1326 2614
rect 1266 2514 1326 2574
rect 1266 2474 1276 2514
rect 1316 2474 1326 2514
rect 1266 2458 1326 2474
rect 1410 2614 1470 2630
rect 1410 2574 1420 2614
rect 1460 2574 1470 2614
rect 1410 2514 1470 2574
rect 1410 2474 1420 2514
rect 1460 2474 1470 2514
rect 1410 2458 1470 2474
rect 1554 2614 1614 2630
rect 1554 2574 1564 2614
rect 1604 2574 1614 2614
rect 1554 2514 1614 2574
rect 1554 2474 1564 2514
rect 1604 2474 1614 2514
rect 1554 2458 1614 2474
rect 1842 2614 1902 2630
rect 1842 2574 1852 2614
rect 1892 2574 1902 2614
rect 1842 2514 1902 2574
rect 1842 2474 1852 2514
rect 1892 2474 1902 2514
rect 1842 2458 1902 2474
rect 1986 2614 2046 2630
rect 1986 2574 1996 2614
rect 2036 2574 2046 2614
rect 1986 2514 2046 2574
rect 1986 2474 1996 2514
rect 2036 2474 2046 2514
rect 1986 2458 2046 2474
rect 2130 2614 2190 2630
rect 2130 2574 2140 2614
rect 2180 2574 2190 2614
rect 2130 2514 2190 2574
rect 2130 2474 2140 2514
rect 2180 2474 2190 2514
rect 2130 2458 2190 2474
rect 2418 2614 2478 2630
rect 2418 2574 2428 2614
rect 2468 2574 2478 2614
rect 2418 2514 2478 2574
rect 2418 2474 2428 2514
rect 2468 2474 2478 2514
rect 2418 2458 2478 2474
rect 2562 2614 2622 2630
rect 2562 2574 2572 2614
rect 2612 2574 2622 2614
rect 2562 2514 2622 2574
rect 2562 2474 2572 2514
rect 2612 2474 2622 2514
rect 2562 2458 2622 2474
rect 2706 2614 2766 2630
rect 2706 2574 2716 2614
rect 2756 2574 2766 2614
rect 2706 2514 2766 2574
rect 2706 2474 2716 2514
rect 2756 2474 2766 2514
rect 2706 2458 2766 2474
rect 2994 2614 3054 2630
rect 2994 2574 3004 2614
rect 3044 2574 3054 2614
rect 2994 2514 3054 2574
rect 2994 2474 3004 2514
rect 3044 2474 3054 2514
rect 2994 2458 3054 2474
rect 3138 2614 3198 2630
rect 3138 2574 3148 2614
rect 3188 2574 3198 2614
rect 3138 2514 3198 2574
rect 3138 2474 3148 2514
rect 3188 2474 3198 2514
rect 3138 2458 3198 2474
rect 3282 2614 3342 2630
rect 3282 2574 3292 2614
rect 3332 2574 3342 2614
rect 3282 2514 3342 2574
rect 3282 2474 3292 2514
rect 3332 2474 3342 2514
rect 3282 2458 3342 2474
rect 3570 2588 3630 2630
rect 3570 2500 3580 2588
rect 3620 2500 3630 2588
rect 3570 2458 3630 2500
rect 3714 2588 3774 2630
rect 3714 2500 3724 2588
rect 3764 2500 3774 2588
rect 3714 2458 3774 2500
rect 3858 2588 3918 2630
rect 3858 2500 3868 2588
rect 3908 2500 3918 2588
rect 3858 2458 3918 2500
rect 4146 2614 4206 2630
rect 4146 2574 4156 2614
rect 4196 2574 4206 2614
rect 4146 2514 4206 2574
rect 4146 2474 4156 2514
rect 4196 2474 4206 2514
rect 4146 2458 4206 2474
rect 4290 2614 4350 2630
rect 4290 2574 4300 2614
rect 4340 2574 4350 2614
rect 4290 2514 4350 2574
rect 4290 2474 4300 2514
rect 4340 2474 4350 2514
rect 4290 2458 4350 2474
rect 4434 2614 4494 2630
rect 4434 2574 4444 2614
rect 4484 2574 4494 2614
rect 4434 2514 4494 2574
rect 4434 2474 4444 2514
rect 4484 2474 4494 2514
rect 4434 2458 4494 2474
rect 4722 2614 4782 2630
rect 4722 2574 4732 2614
rect 4772 2574 4782 2614
rect 4722 2514 4782 2574
rect 4722 2474 4732 2514
rect 4772 2474 4782 2514
rect 4722 2458 4782 2474
rect 4866 2614 4926 2630
rect 4866 2574 4876 2614
rect 4916 2574 4926 2614
rect 4866 2514 4926 2574
rect 4866 2474 4876 2514
rect 4916 2474 4926 2514
rect 4866 2458 4926 2474
rect 5010 2614 5070 2630
rect 5010 2574 5020 2614
rect 5060 2574 5070 2614
rect 5010 2514 5070 2574
rect 5010 2474 5020 2514
rect 5060 2474 5070 2514
rect 5010 2458 5070 2474
rect 5298 2614 5358 2630
rect 5298 2574 5308 2614
rect 5348 2574 5358 2614
rect 5298 2514 5358 2574
rect 5298 2474 5308 2514
rect 5348 2474 5358 2514
rect 5298 2458 5358 2474
rect 5442 2614 5502 2630
rect 5442 2574 5452 2614
rect 5492 2574 5502 2614
rect 5442 2514 5502 2574
rect 5442 2474 5452 2514
rect 5492 2474 5502 2514
rect 5442 2458 5502 2474
rect 5586 2614 5646 2630
rect 5586 2574 5596 2614
rect 5636 2574 5646 2614
rect 5586 2514 5646 2574
rect 5586 2474 5596 2514
rect 5636 2474 5646 2514
rect 5586 2458 5646 2474
rect 5874 2614 5934 2630
rect 5874 2574 5884 2614
rect 5924 2574 5934 2614
rect 5874 2514 5934 2574
rect 5874 2474 5884 2514
rect 5924 2474 5934 2514
rect 5874 2458 5934 2474
rect 6018 2614 6078 2630
rect 6018 2574 6028 2614
rect 6068 2574 6078 2614
rect 6018 2514 6078 2574
rect 6018 2474 6028 2514
rect 6068 2474 6078 2514
rect 6018 2458 6078 2474
rect 6162 2614 6222 2630
rect 6162 2574 6172 2614
rect 6212 2574 6222 2614
rect 6162 2514 6222 2574
rect 6162 2474 6172 2514
rect 6212 2474 6222 2514
rect 6162 2458 6222 2474
rect 6450 2614 6510 2630
rect 6450 2574 6460 2614
rect 6500 2574 6510 2614
rect 6450 2514 6510 2574
rect 6450 2474 6460 2514
rect 6500 2474 6510 2514
rect 6450 2458 6510 2474
rect 6594 2614 6654 2630
rect 6594 2574 6604 2614
rect 6644 2574 6654 2614
rect 6594 2514 6654 2574
rect 6594 2474 6604 2514
rect 6644 2474 6654 2514
rect 6594 2458 6654 2474
rect 6738 2614 6798 2630
rect 6738 2574 6748 2614
rect 6788 2574 6798 2614
rect 6738 2514 6798 2574
rect 6738 2474 6748 2514
rect 6788 2474 6798 2514
rect 6738 2458 6798 2474
rect 7026 2588 7086 2630
rect 7026 2500 7036 2588
rect 7076 2500 7086 2588
rect 7026 2458 7086 2500
rect 7170 2588 7230 2630
rect 7170 2500 7180 2588
rect 7220 2500 7230 2588
rect 7170 2458 7230 2500
rect 7314 2588 7374 2630
rect 7314 2500 7324 2588
rect 7364 2500 7374 2588
rect 7314 2458 7374 2500
rect 7602 2614 7662 2630
rect 7602 2574 7612 2614
rect 7652 2574 7662 2614
rect 7602 2514 7662 2574
rect 7602 2474 7612 2514
rect 7652 2474 7662 2514
rect 7602 2458 7662 2474
rect 7746 2614 7806 2630
rect 7746 2574 7756 2614
rect 7796 2574 7806 2614
rect 7746 2514 7806 2574
rect 7746 2474 7756 2514
rect 7796 2474 7806 2514
rect 7746 2458 7806 2474
rect 7890 2614 7950 2630
rect 7890 2574 7900 2614
rect 7940 2574 7950 2614
rect 7890 2514 7950 2574
rect 7890 2474 7900 2514
rect 7940 2474 7950 2514
rect 7890 2458 7950 2474
rect 8178 2614 8238 2630
rect 8178 2574 8188 2614
rect 8228 2574 8238 2614
rect 8178 2514 8238 2574
rect 8178 2474 8188 2514
rect 8228 2474 8238 2514
rect 8178 2458 8238 2474
rect 8322 2614 8382 2630
rect 8322 2574 8332 2614
rect 8372 2574 8382 2614
rect 8322 2514 8382 2574
rect 8322 2474 8332 2514
rect 8372 2474 8382 2514
rect 8322 2458 8382 2474
rect 8466 2614 8526 2630
rect 8466 2574 8476 2614
rect 8516 2574 8526 2614
rect 8466 2514 8526 2574
rect 8466 2474 8476 2514
rect 8516 2474 8526 2514
rect 8466 2458 8526 2474
rect 8754 2614 8814 2630
rect 8754 2574 8764 2614
rect 8804 2574 8814 2614
rect 8754 2514 8814 2574
rect 8754 2474 8764 2514
rect 8804 2474 8814 2514
rect 8754 2458 8814 2474
rect 8898 2614 8958 2630
rect 8898 2574 8908 2614
rect 8948 2574 8958 2614
rect 8898 2514 8958 2574
rect 8898 2474 8908 2514
rect 8948 2474 8958 2514
rect 8898 2458 8958 2474
rect 9042 2614 9102 2630
rect 9042 2574 9052 2614
rect 9092 2574 9102 2614
rect 9042 2514 9102 2574
rect 9042 2474 9052 2514
rect 9092 2474 9102 2514
rect 9042 2458 9102 2474
rect 9330 2614 9390 2630
rect 9330 2574 9340 2614
rect 9380 2574 9390 2614
rect 9330 2514 9390 2574
rect 9330 2474 9340 2514
rect 9380 2474 9390 2514
rect 9330 2458 9390 2474
rect 9474 2614 9534 2630
rect 9474 2574 9484 2614
rect 9524 2574 9534 2614
rect 9474 2514 9534 2574
rect 9474 2474 9484 2514
rect 9524 2474 9534 2514
rect 9474 2458 9534 2474
rect 9618 2614 9678 2630
rect 9618 2574 9628 2614
rect 9668 2574 9678 2614
rect 9618 2514 9678 2574
rect 9618 2474 9628 2514
rect 9668 2474 9678 2514
rect 9618 2458 9678 2474
rect 10194 2614 10254 2630
rect 10194 2574 10204 2614
rect 10244 2574 10254 2614
rect 10194 2514 10254 2574
rect 10194 2474 10204 2514
rect 10244 2474 10254 2514
rect 10194 2458 10254 2474
rect 10338 2614 10398 2630
rect 10338 2574 10348 2614
rect 10388 2574 10398 2614
rect 10338 2514 10398 2574
rect 10338 2474 10348 2514
rect 10388 2474 10398 2514
rect 10338 2458 10398 2474
rect 10482 2614 10542 2630
rect 10482 2574 10492 2614
rect 10532 2574 10542 2614
rect 10482 2514 10542 2574
rect 10482 2474 10492 2514
rect 10532 2474 10542 2514
rect 10482 2458 10542 2474
rect 10770 2614 10830 2630
rect 10770 2574 10780 2614
rect 10820 2574 10830 2614
rect 10770 2514 10830 2574
rect 10770 2474 10780 2514
rect 10820 2474 10830 2514
rect 10770 2458 10830 2474
rect 10914 2614 10974 2630
rect 10914 2574 10924 2614
rect 10964 2574 10974 2614
rect 10914 2514 10974 2574
rect 10914 2474 10924 2514
rect 10964 2474 10974 2514
rect 10914 2458 10974 2474
rect 11058 2614 11118 2630
rect 11058 2574 11068 2614
rect 11108 2574 11118 2614
rect 11058 2514 11118 2574
rect 11058 2474 11068 2514
rect 11108 2474 11118 2514
rect 11058 2458 11118 2474
rect 11346 2588 11406 2630
rect 11346 2500 11356 2588
rect 11396 2500 11406 2588
rect 11346 2458 11406 2500
rect 11490 2588 11550 2630
rect 11490 2500 11500 2588
rect 11540 2500 11550 2588
rect 11490 2458 11550 2500
rect 11634 2588 11694 2630
rect 11634 2500 11644 2588
rect 11684 2500 11694 2588
rect 11634 2458 11694 2500
rect 11922 2614 11982 2630
rect 11922 2574 11932 2614
rect 11972 2574 11982 2614
rect 11922 2514 11982 2574
rect 11922 2474 11932 2514
rect 11972 2474 11982 2514
rect 11922 2458 11982 2474
rect 12066 2614 12126 2630
rect 12066 2574 12076 2614
rect 12116 2574 12126 2614
rect 12066 2514 12126 2574
rect 12066 2474 12076 2514
rect 12116 2474 12126 2514
rect 12066 2458 12126 2474
rect 12210 2614 12270 2630
rect 12210 2574 12220 2614
rect 12260 2574 12270 2614
rect 12210 2514 12270 2574
rect 12210 2474 12220 2514
rect 12260 2474 12270 2514
rect 12210 2458 12270 2474
rect 12498 2614 12558 2630
rect 12498 2574 12508 2614
rect 12548 2574 12558 2614
rect 12498 2514 12558 2574
rect 12498 2474 12508 2514
rect 12548 2474 12558 2514
rect 12498 2458 12558 2474
rect 12642 2614 12702 2630
rect 12642 2574 12652 2614
rect 12692 2574 12702 2614
rect 12642 2514 12702 2574
rect 12642 2474 12652 2514
rect 12692 2474 12702 2514
rect 12642 2458 12702 2474
rect 12786 2614 12846 2630
rect 12786 2574 12796 2614
rect 12836 2574 12846 2614
rect 12786 2514 12846 2574
rect 12786 2474 12796 2514
rect 12836 2474 12846 2514
rect 12786 2458 12846 2474
rect 13650 2614 13710 2630
rect 13650 2574 13660 2614
rect 13700 2574 13710 2614
rect 13650 2514 13710 2574
rect 13650 2474 13660 2514
rect 13700 2474 13710 2514
rect 13650 2458 13710 2474
rect 13794 2614 13854 2630
rect 13794 2574 13804 2614
rect 13844 2574 13854 2614
rect 13794 2514 13854 2574
rect 13794 2474 13804 2514
rect 13844 2474 13854 2514
rect 13794 2458 13854 2474
rect 13938 2614 13998 2630
rect 13938 2574 13948 2614
rect 13988 2574 13998 2614
rect 13938 2514 13998 2574
rect 13938 2474 13948 2514
rect 13988 2474 13998 2514
rect 13938 2458 13998 2474
rect 14226 2614 14286 2630
rect 14226 2574 14236 2614
rect 14276 2574 14286 2614
rect 14226 2514 14286 2574
rect 14226 2474 14236 2514
rect 14276 2474 14286 2514
rect 14226 2458 14286 2474
rect 14370 2614 14430 2630
rect 14370 2574 14380 2614
rect 14420 2574 14430 2614
rect 14370 2514 14430 2574
rect 14370 2474 14380 2514
rect 14420 2474 14430 2514
rect 14370 2458 14430 2474
rect 14514 2614 14574 2630
rect 14514 2574 14524 2614
rect 14564 2574 14574 2614
rect 14514 2514 14574 2574
rect 14514 2474 14524 2514
rect 14564 2474 14574 2514
rect 14514 2458 14574 2474
rect 14802 2614 14862 2630
rect 14802 2574 14812 2614
rect 14852 2574 14862 2614
rect 14802 2514 14862 2574
rect 14802 2474 14812 2514
rect 14852 2474 14862 2514
rect 14802 2458 14862 2474
rect 14946 2614 15006 2630
rect 14946 2574 14956 2614
rect 14996 2574 15006 2614
rect 14946 2514 15006 2574
rect 14946 2474 14956 2514
rect 14996 2474 15006 2514
rect 14946 2458 15006 2474
rect 15090 2614 15150 2630
rect 15090 2574 15100 2614
rect 15140 2574 15150 2614
rect 15090 2514 15150 2574
rect 15090 2474 15100 2514
rect 15140 2474 15150 2514
rect 15090 2458 15150 2474
rect 15378 2588 15438 2630
rect 15378 2500 15388 2588
rect 15428 2500 15438 2588
rect 15378 2458 15438 2500
rect 15522 2588 15582 2630
rect 15522 2500 15532 2588
rect 15572 2500 15582 2588
rect 15522 2458 15582 2500
rect 15666 2588 15726 2630
rect 15666 2500 15676 2588
rect 15716 2500 15726 2588
rect 15666 2458 15726 2500
rect 15954 2588 16014 2630
rect 15954 2500 15964 2588
rect 16004 2500 16014 2588
rect 15954 2458 16014 2500
rect 16098 2588 16158 2630
rect 16098 2500 16108 2588
rect 16148 2500 16158 2588
rect 16098 2458 16158 2500
rect 16242 2588 16302 2630
rect 16242 2500 16252 2588
rect 16292 2500 16302 2588
rect 16242 2458 16302 2500
rect 16530 2614 16590 2630
rect 16530 2574 16540 2614
rect 16580 2574 16590 2614
rect 16530 2514 16590 2574
rect 16530 2474 16540 2514
rect 16580 2474 16590 2514
rect 16530 2458 16590 2474
rect 16674 2614 16734 2630
rect 16674 2574 16684 2614
rect 16724 2574 16734 2614
rect 16674 2514 16734 2574
rect 16674 2474 16684 2514
rect 16724 2474 16734 2514
rect 16674 2458 16734 2474
rect 16818 2614 16878 2630
rect 16818 2574 16828 2614
rect 16868 2574 16878 2614
rect 16818 2514 16878 2574
rect 16818 2474 16828 2514
rect 16868 2474 16878 2514
rect 16818 2458 16878 2474
rect 16962 2614 17022 2630
rect 16962 2574 16972 2614
rect 17012 2574 17022 2614
rect 16962 2514 17022 2574
rect 16962 2474 16972 2514
rect 17012 2474 17022 2514
rect 16962 2458 17022 2474
rect 17106 2614 17166 2630
rect 17106 2574 17116 2614
rect 17156 2574 17166 2614
rect 17106 2514 17166 2574
rect 17106 2474 17116 2514
rect 17156 2474 17166 2514
rect 17106 2458 17166 2474
rect 17250 2614 17310 2630
rect 17250 2574 17260 2614
rect 17300 2574 17310 2614
rect 17250 2514 17310 2574
rect 17250 2474 17260 2514
rect 17300 2474 17310 2514
rect 17250 2458 17310 2474
rect 17394 2614 17454 2630
rect 17394 2574 17404 2614
rect 17444 2574 17454 2614
rect 17394 2514 17454 2574
rect 17394 2474 17404 2514
rect 17444 2474 17454 2514
rect 17394 2458 17454 2474
rect 17538 2614 17598 2630
rect 17538 2574 17548 2614
rect 17588 2574 17598 2614
rect 17538 2514 17598 2574
rect 17538 2474 17548 2514
rect 17588 2474 17598 2514
rect 17538 2458 17598 2474
rect 17682 2614 17742 2630
rect 17682 2574 17692 2614
rect 17732 2574 17742 2614
rect 17682 2514 17742 2574
rect 17682 2474 17692 2514
rect 17732 2474 17742 2514
rect 17682 2458 17742 2474
rect 17826 2614 17886 2630
rect 17826 2574 17836 2614
rect 17876 2574 17886 2614
rect 17826 2514 17886 2574
rect 17826 2474 17836 2514
rect 17876 2474 17886 2514
rect 17826 2458 17886 2474
rect 17970 2614 18030 2630
rect 17970 2574 17980 2614
rect 18020 2574 18030 2614
rect 17970 2514 18030 2574
rect 17970 2474 17980 2514
rect 18020 2474 18030 2514
rect 17970 2458 18030 2474
rect 18114 2614 18174 2630
rect 18114 2574 18124 2614
rect 18164 2574 18174 2614
rect 18114 2514 18174 2574
rect 18114 2474 18124 2514
rect 18164 2474 18174 2514
rect 18114 2458 18174 2474
rect 18258 2614 18318 2630
rect 18258 2574 18268 2614
rect 18308 2574 18318 2614
rect 18258 2514 18318 2574
rect 18258 2474 18268 2514
rect 18308 2474 18318 2514
rect 18258 2458 18318 2474
rect 18402 2614 18462 2630
rect 18402 2574 18412 2614
rect 18452 2574 18462 2614
rect 18402 2514 18462 2574
rect 18402 2474 18412 2514
rect 18452 2474 18462 2514
rect 18402 2458 18462 2474
rect 18546 2614 18606 2630
rect 18546 2574 18556 2614
rect 18596 2574 18606 2614
rect 18546 2514 18606 2574
rect 18546 2474 18556 2514
rect 18596 2474 18606 2514
rect 18546 2458 18606 2474
rect 18690 2614 18750 2630
rect 18690 2574 18700 2614
rect 18740 2574 18750 2614
rect 18690 2514 18750 2574
rect 18690 2474 18700 2514
rect 18740 2474 18750 2514
rect 18690 2458 18750 2474
rect 18834 2614 18894 2630
rect 18834 2574 18844 2614
rect 18884 2574 18894 2614
rect 18834 2514 18894 2574
rect 18834 2474 18844 2514
rect 18884 2474 18894 2514
rect 18834 2458 18894 2474
rect 18978 2614 19038 2630
rect 18978 2574 18988 2614
rect 19028 2574 19038 2614
rect 18978 2514 19038 2574
rect 18978 2474 18988 2514
rect 19028 2474 19038 2514
rect 18978 2458 19038 2474
rect 19122 2614 19182 2630
rect 19122 2574 19132 2614
rect 19172 2574 19182 2614
rect 19122 2514 19182 2574
rect 19122 2474 19132 2514
rect 19172 2474 19182 2514
rect 19122 2458 19182 2474
rect 19266 2614 19326 2630
rect 19266 2574 19276 2614
rect 19316 2574 19326 2614
rect 19266 2514 19326 2574
rect 19266 2474 19276 2514
rect 19316 2474 19326 2514
rect 19266 2458 19326 2474
rect 19410 2614 19470 2630
rect 19410 2574 19420 2614
rect 19460 2574 19470 2614
rect 19410 2514 19470 2574
rect 19410 2474 19420 2514
rect 19460 2474 19470 2514
rect 19410 2458 19470 2474
rect 19554 2614 19614 2630
rect 19554 2574 19564 2614
rect 19604 2574 19614 2614
rect 19554 2514 19614 2574
rect 19554 2474 19564 2514
rect 19604 2474 19614 2514
rect 19554 2458 19614 2474
rect 19698 2614 19758 2630
rect 19698 2574 19708 2614
rect 19748 2574 19758 2614
rect 19698 2514 19758 2574
rect 19698 2474 19708 2514
rect 19748 2474 19758 2514
rect 19698 2458 19758 2474
rect 19842 2614 19902 2630
rect 19842 2574 19852 2614
rect 19892 2574 19902 2614
rect 19842 2514 19902 2574
rect 19842 2474 19852 2514
rect 19892 2474 19902 2514
rect 19842 2458 19902 2474
rect 19986 2614 20046 2630
rect 19986 2574 19996 2614
rect 20036 2574 20046 2614
rect 19986 2514 20046 2574
rect 19986 2474 19996 2514
rect 20036 2474 20046 2514
rect 19986 2458 20046 2474
rect 114 1532 174 1574
rect 114 1444 124 1532
rect 164 1444 174 1532
rect 114 1402 174 1444
rect 258 1532 318 1574
rect 258 1444 268 1532
rect 308 1444 318 1532
rect 258 1402 318 1444
rect 402 1532 462 1574
rect 402 1444 412 1532
rect 452 1444 462 1532
rect 402 1402 462 1444
rect 690 1558 750 1574
rect 690 1518 700 1558
rect 740 1518 750 1558
rect 690 1458 750 1518
rect 690 1418 700 1458
rect 740 1418 750 1458
rect 690 1402 750 1418
rect 834 1558 894 1574
rect 834 1518 844 1558
rect 884 1518 894 1558
rect 834 1458 894 1518
rect 834 1418 844 1458
rect 884 1418 894 1458
rect 834 1402 894 1418
rect 978 1558 1038 1574
rect 978 1518 988 1558
rect 1028 1518 1038 1558
rect 978 1458 1038 1518
rect 978 1418 988 1458
rect 1028 1418 1038 1458
rect 978 1402 1038 1418
rect 1266 1558 1326 1574
rect 1266 1518 1276 1558
rect 1316 1518 1326 1558
rect 1266 1458 1326 1518
rect 1266 1418 1276 1458
rect 1316 1418 1326 1458
rect 1266 1402 1326 1418
rect 1410 1558 1470 1574
rect 1410 1518 1420 1558
rect 1460 1518 1470 1558
rect 1410 1458 1470 1518
rect 1410 1418 1420 1458
rect 1460 1418 1470 1458
rect 1410 1402 1470 1418
rect 1554 1558 1614 1574
rect 1554 1518 1564 1558
rect 1604 1518 1614 1558
rect 1554 1458 1614 1518
rect 1554 1418 1564 1458
rect 1604 1418 1614 1458
rect 1554 1402 1614 1418
rect 1842 1558 1902 1574
rect 1842 1518 1852 1558
rect 1892 1518 1902 1558
rect 1842 1458 1902 1518
rect 1842 1418 1852 1458
rect 1892 1418 1902 1458
rect 1842 1402 1902 1418
rect 1986 1558 2046 1574
rect 1986 1518 1996 1558
rect 2036 1518 2046 1558
rect 1986 1458 2046 1518
rect 1986 1418 1996 1458
rect 2036 1418 2046 1458
rect 1986 1402 2046 1418
rect 2130 1558 2190 1574
rect 2130 1518 2140 1558
rect 2180 1518 2190 1558
rect 2130 1458 2190 1518
rect 2130 1418 2140 1458
rect 2180 1418 2190 1458
rect 2130 1402 2190 1418
rect 2994 1558 3054 1574
rect 2994 1518 3004 1558
rect 3044 1518 3054 1558
rect 2994 1458 3054 1518
rect 2994 1418 3004 1458
rect 3044 1418 3054 1458
rect 2994 1402 3054 1418
rect 3138 1558 3198 1574
rect 3138 1518 3148 1558
rect 3188 1518 3198 1558
rect 3138 1458 3198 1518
rect 3138 1418 3148 1458
rect 3188 1418 3198 1458
rect 3138 1402 3198 1418
rect 3282 1558 3342 1574
rect 3282 1518 3292 1558
rect 3332 1518 3342 1558
rect 3282 1458 3342 1518
rect 3282 1418 3292 1458
rect 3332 1418 3342 1458
rect 3282 1402 3342 1418
rect 3570 1558 3630 1574
rect 3570 1518 3580 1558
rect 3620 1518 3630 1558
rect 3570 1458 3630 1518
rect 3570 1418 3580 1458
rect 3620 1418 3630 1458
rect 3570 1402 3630 1418
rect 3714 1558 3774 1574
rect 3714 1518 3724 1558
rect 3764 1518 3774 1558
rect 3714 1458 3774 1518
rect 3714 1418 3724 1458
rect 3764 1418 3774 1458
rect 3714 1402 3774 1418
rect 3858 1558 3918 1574
rect 3858 1518 3868 1558
rect 3908 1518 3918 1558
rect 3858 1458 3918 1518
rect 3858 1418 3868 1458
rect 3908 1418 3918 1458
rect 3858 1402 3918 1418
rect 4146 1558 4206 1574
rect 4146 1518 4156 1558
rect 4196 1518 4206 1558
rect 4146 1458 4206 1518
rect 4146 1418 4156 1458
rect 4196 1418 4206 1458
rect 4146 1402 4206 1418
rect 4290 1558 4350 1574
rect 4290 1518 4300 1558
rect 4340 1518 4350 1558
rect 4290 1458 4350 1518
rect 4290 1418 4300 1458
rect 4340 1418 4350 1458
rect 4290 1402 4350 1418
rect 4434 1558 4494 1574
rect 4434 1518 4444 1558
rect 4484 1518 4494 1558
rect 4434 1458 4494 1518
rect 4434 1418 4444 1458
rect 4484 1418 4494 1458
rect 4434 1402 4494 1418
rect 4722 1532 4782 1574
rect 4722 1444 4732 1532
rect 4772 1444 4782 1532
rect 4722 1402 4782 1444
rect 4866 1532 4926 1574
rect 4866 1444 4876 1532
rect 4916 1444 4926 1532
rect 4866 1402 4926 1444
rect 5010 1532 5070 1574
rect 5010 1444 5020 1532
rect 5060 1444 5070 1532
rect 5010 1402 5070 1444
rect 5298 1532 5358 1574
rect 5298 1444 5308 1532
rect 5348 1444 5358 1532
rect 5298 1402 5358 1444
rect 5442 1532 5502 1574
rect 5442 1444 5452 1532
rect 5492 1444 5502 1532
rect 5442 1402 5502 1444
rect 5586 1532 5646 1574
rect 5586 1444 5596 1532
rect 5636 1444 5646 1532
rect 5586 1402 5646 1444
rect 5874 1558 5934 1574
rect 5874 1518 5884 1558
rect 5924 1518 5934 1558
rect 5874 1458 5934 1518
rect 5874 1418 5884 1458
rect 5924 1418 5934 1458
rect 5874 1402 5934 1418
rect 6018 1558 6078 1574
rect 6018 1518 6028 1558
rect 6068 1518 6078 1558
rect 6018 1458 6078 1518
rect 6018 1418 6028 1458
rect 6068 1418 6078 1458
rect 6018 1402 6078 1418
rect 6162 1558 6222 1574
rect 6162 1518 6172 1558
rect 6212 1518 6222 1558
rect 6162 1458 6222 1518
rect 6162 1418 6172 1458
rect 6212 1418 6222 1458
rect 6162 1402 6222 1418
rect 6450 1558 6510 1574
rect 6450 1518 6460 1558
rect 6500 1518 6510 1558
rect 6450 1458 6510 1518
rect 6450 1418 6460 1458
rect 6500 1418 6510 1458
rect 6450 1402 6510 1418
rect 6594 1558 6654 1574
rect 6594 1518 6604 1558
rect 6644 1518 6654 1558
rect 6594 1458 6654 1518
rect 6594 1418 6604 1458
rect 6644 1418 6654 1458
rect 6594 1402 6654 1418
rect 6738 1558 6798 1574
rect 6738 1518 6748 1558
rect 6788 1518 6798 1558
rect 6738 1458 6798 1518
rect 6738 1418 6748 1458
rect 6788 1418 6798 1458
rect 6738 1402 6798 1418
rect 7026 1558 7086 1574
rect 7026 1518 7036 1558
rect 7076 1518 7086 1558
rect 7026 1458 7086 1518
rect 7026 1418 7036 1458
rect 7076 1418 7086 1458
rect 7026 1402 7086 1418
rect 7170 1558 7230 1574
rect 7170 1518 7180 1558
rect 7220 1518 7230 1558
rect 7170 1458 7230 1518
rect 7170 1418 7180 1458
rect 7220 1418 7230 1458
rect 7170 1402 7230 1418
rect 7314 1558 7374 1574
rect 7314 1518 7324 1558
rect 7364 1518 7374 1558
rect 7314 1458 7374 1518
rect 7314 1418 7324 1458
rect 7364 1418 7374 1458
rect 7314 1402 7374 1418
rect 7602 1558 7662 1574
rect 7602 1518 7612 1558
rect 7652 1518 7662 1558
rect 7602 1458 7662 1518
rect 7602 1418 7612 1458
rect 7652 1418 7662 1458
rect 7602 1402 7662 1418
rect 7746 1558 7806 1574
rect 7746 1518 7756 1558
rect 7796 1518 7806 1558
rect 7746 1458 7806 1518
rect 7746 1418 7756 1458
rect 7796 1418 7806 1458
rect 7746 1402 7806 1418
rect 7890 1558 7950 1574
rect 7890 1518 7900 1558
rect 7940 1518 7950 1558
rect 7890 1458 7950 1518
rect 7890 1418 7900 1458
rect 7940 1418 7950 1458
rect 7890 1402 7950 1418
rect 8178 1558 8238 1574
rect 8178 1518 8188 1558
rect 8228 1518 8238 1558
rect 8178 1458 8238 1518
rect 8178 1418 8188 1458
rect 8228 1418 8238 1458
rect 8178 1402 8238 1418
rect 8322 1558 8382 1574
rect 8322 1518 8332 1558
rect 8372 1518 8382 1558
rect 8322 1458 8382 1518
rect 8322 1418 8332 1458
rect 8372 1418 8382 1458
rect 8322 1402 8382 1418
rect 8466 1558 8526 1574
rect 8466 1518 8476 1558
rect 8516 1518 8526 1558
rect 8466 1458 8526 1518
rect 8466 1418 8476 1458
rect 8516 1418 8526 1458
rect 8466 1402 8526 1418
rect 8754 1532 8814 1574
rect 8754 1444 8764 1532
rect 8804 1444 8814 1532
rect 8754 1402 8814 1444
rect 8898 1532 8958 1574
rect 8898 1444 8908 1532
rect 8948 1444 8958 1532
rect 8898 1402 8958 1444
rect 9042 1532 9102 1574
rect 9042 1444 9052 1532
rect 9092 1444 9102 1532
rect 9042 1402 9102 1444
rect 9330 1558 9390 1574
rect 9330 1518 9340 1558
rect 9380 1518 9390 1558
rect 9330 1458 9390 1518
rect 9330 1418 9340 1458
rect 9380 1418 9390 1458
rect 9330 1402 9390 1418
rect 9474 1558 9534 1574
rect 9474 1518 9484 1558
rect 9524 1518 9534 1558
rect 9474 1458 9534 1518
rect 9474 1418 9484 1458
rect 9524 1418 9534 1458
rect 9474 1402 9534 1418
rect 9618 1558 9678 1574
rect 9618 1518 9628 1558
rect 9668 1518 9678 1558
rect 9618 1458 9678 1518
rect 9618 1418 9628 1458
rect 9668 1418 9678 1458
rect 9618 1402 9678 1418
rect 9906 1558 9966 1574
rect 9906 1518 9916 1558
rect 9956 1518 9966 1558
rect 9906 1458 9966 1518
rect 9906 1418 9916 1458
rect 9956 1418 9966 1458
rect 9906 1402 9966 1418
rect 10050 1558 10110 1574
rect 10050 1518 10060 1558
rect 10100 1518 10110 1558
rect 10050 1458 10110 1518
rect 10050 1418 10060 1458
rect 10100 1418 10110 1458
rect 10050 1402 10110 1418
rect 10194 1558 10254 1574
rect 10194 1518 10204 1558
rect 10244 1518 10254 1558
rect 10194 1458 10254 1518
rect 10194 1418 10204 1458
rect 10244 1418 10254 1458
rect 10194 1402 10254 1418
rect 10482 1558 10542 1574
rect 10482 1518 10492 1558
rect 10532 1518 10542 1558
rect 10482 1458 10542 1518
rect 10482 1418 10492 1458
rect 10532 1418 10542 1458
rect 10482 1402 10542 1418
rect 10626 1558 10686 1574
rect 10626 1518 10636 1558
rect 10676 1518 10686 1558
rect 10626 1458 10686 1518
rect 10626 1418 10636 1458
rect 10676 1418 10686 1458
rect 10626 1402 10686 1418
rect 10770 1558 10830 1574
rect 10770 1518 10780 1558
rect 10820 1518 10830 1558
rect 10770 1458 10830 1518
rect 10770 1418 10780 1458
rect 10820 1418 10830 1458
rect 10770 1402 10830 1418
rect 11058 1558 11118 1574
rect 11058 1518 11068 1558
rect 11108 1518 11118 1558
rect 11058 1458 11118 1518
rect 11058 1418 11068 1458
rect 11108 1418 11118 1458
rect 11058 1402 11118 1418
rect 11202 1558 11262 1574
rect 11202 1518 11212 1558
rect 11252 1518 11262 1558
rect 11202 1458 11262 1518
rect 11202 1418 11212 1458
rect 11252 1418 11262 1458
rect 11202 1402 11262 1418
rect 11346 1558 11406 1574
rect 11346 1518 11356 1558
rect 11396 1518 11406 1558
rect 11346 1458 11406 1518
rect 11346 1418 11356 1458
rect 11396 1418 11406 1458
rect 11346 1402 11406 1418
rect 11922 1558 11982 1574
rect 11922 1518 11932 1558
rect 11972 1518 11982 1558
rect 11922 1458 11982 1518
rect 11922 1418 11932 1458
rect 11972 1418 11982 1458
rect 11922 1402 11982 1418
rect 12066 1558 12126 1574
rect 12066 1518 12076 1558
rect 12116 1518 12126 1558
rect 12066 1458 12126 1518
rect 12066 1418 12076 1458
rect 12116 1418 12126 1458
rect 12066 1402 12126 1418
rect 12210 1558 12270 1574
rect 12210 1518 12220 1558
rect 12260 1518 12270 1558
rect 12210 1458 12270 1518
rect 12210 1418 12220 1458
rect 12260 1418 12270 1458
rect 12210 1402 12270 1418
rect 12498 1558 12558 1574
rect 12498 1518 12508 1558
rect 12548 1518 12558 1558
rect 12498 1458 12558 1518
rect 12498 1418 12508 1458
rect 12548 1418 12558 1458
rect 12498 1402 12558 1418
rect 12642 1558 12702 1574
rect 12642 1518 12652 1558
rect 12692 1518 12702 1558
rect 12642 1458 12702 1518
rect 12642 1418 12652 1458
rect 12692 1418 12702 1458
rect 12642 1402 12702 1418
rect 12786 1558 12846 1574
rect 12786 1518 12796 1558
rect 12836 1518 12846 1558
rect 12786 1458 12846 1518
rect 12786 1418 12796 1458
rect 12836 1418 12846 1458
rect 12786 1402 12846 1418
rect 13074 1558 13134 1574
rect 13074 1518 13084 1558
rect 13124 1518 13134 1558
rect 13074 1458 13134 1518
rect 13074 1418 13084 1458
rect 13124 1418 13134 1458
rect 13074 1402 13134 1418
rect 13218 1558 13278 1574
rect 13218 1518 13228 1558
rect 13268 1518 13278 1558
rect 13218 1458 13278 1518
rect 13218 1418 13228 1458
rect 13268 1418 13278 1458
rect 13218 1402 13278 1418
rect 13362 1558 13422 1574
rect 13362 1518 13372 1558
rect 13412 1518 13422 1558
rect 13362 1458 13422 1518
rect 13362 1418 13372 1458
rect 13412 1418 13422 1458
rect 13362 1402 13422 1418
rect 13650 1558 13710 1574
rect 13650 1518 13660 1558
rect 13700 1518 13710 1558
rect 13650 1458 13710 1518
rect 13650 1418 13660 1458
rect 13700 1418 13710 1458
rect 13650 1402 13710 1418
rect 13794 1558 13854 1574
rect 13794 1518 13804 1558
rect 13844 1518 13854 1558
rect 13794 1458 13854 1518
rect 13794 1418 13804 1458
rect 13844 1418 13854 1458
rect 13794 1402 13854 1418
rect 13938 1558 13998 1574
rect 13938 1518 13948 1558
rect 13988 1518 13998 1558
rect 13938 1458 13998 1518
rect 13938 1418 13948 1458
rect 13988 1418 13998 1458
rect 13938 1402 13998 1418
rect 14226 1532 14286 1574
rect 14226 1444 14236 1532
rect 14276 1444 14286 1532
rect 14226 1402 14286 1444
rect 14370 1532 14430 1574
rect 14370 1444 14380 1532
rect 14420 1444 14430 1532
rect 14370 1402 14430 1444
rect 14514 1532 14574 1574
rect 14514 1444 14524 1532
rect 14564 1444 14574 1532
rect 14514 1402 14574 1444
rect 14802 1558 14862 1574
rect 14802 1518 14812 1558
rect 14852 1518 14862 1558
rect 14802 1458 14862 1518
rect 14802 1418 14812 1458
rect 14852 1418 14862 1458
rect 14802 1402 14862 1418
rect 14946 1558 15006 1574
rect 14946 1518 14956 1558
rect 14996 1518 15006 1558
rect 14946 1458 15006 1518
rect 14946 1418 14956 1458
rect 14996 1418 15006 1458
rect 14946 1402 15006 1418
rect 15090 1558 15150 1574
rect 15090 1518 15100 1558
rect 15140 1518 15150 1558
rect 15090 1458 15150 1518
rect 15090 1418 15100 1458
rect 15140 1418 15150 1458
rect 15090 1402 15150 1418
rect 15378 1558 15438 1574
rect 15378 1518 15388 1558
rect 15428 1518 15438 1558
rect 15378 1458 15438 1518
rect 15378 1418 15388 1458
rect 15428 1418 15438 1458
rect 15378 1402 15438 1418
rect 15522 1558 15582 1574
rect 15522 1518 15532 1558
rect 15572 1518 15582 1558
rect 15522 1458 15582 1518
rect 15522 1418 15532 1458
rect 15572 1418 15582 1458
rect 15522 1402 15582 1418
rect 15666 1558 15726 1574
rect 15666 1518 15676 1558
rect 15716 1518 15726 1558
rect 15666 1458 15726 1518
rect 15666 1418 15676 1458
rect 15716 1418 15726 1458
rect 15666 1402 15726 1418
rect 15954 1558 16014 1574
rect 15954 1518 15964 1558
rect 16004 1518 16014 1558
rect 15954 1458 16014 1518
rect 15954 1418 15964 1458
rect 16004 1418 16014 1458
rect 15954 1402 16014 1418
rect 16098 1558 16158 1574
rect 16098 1518 16108 1558
rect 16148 1518 16158 1558
rect 16098 1458 16158 1518
rect 16098 1418 16108 1458
rect 16148 1418 16158 1458
rect 16098 1402 16158 1418
rect 16242 1558 16302 1574
rect 16242 1518 16252 1558
rect 16292 1518 16302 1558
rect 16242 1458 16302 1518
rect 16242 1418 16252 1458
rect 16292 1418 16302 1458
rect 16242 1402 16302 1418
rect 16386 1558 16446 1574
rect 16386 1518 16396 1558
rect 16436 1518 16446 1558
rect 16386 1458 16446 1518
rect 16386 1418 16396 1458
rect 16436 1418 16446 1458
rect 16386 1402 16446 1418
rect 16530 1558 16590 1574
rect 16530 1518 16540 1558
rect 16580 1518 16590 1558
rect 16530 1458 16590 1518
rect 16530 1418 16540 1458
rect 16580 1418 16590 1458
rect 16530 1402 16590 1418
rect 16818 1532 16878 1574
rect 16818 1444 16828 1532
rect 16868 1444 16878 1532
rect 16818 1402 16878 1444
rect 16962 1532 17022 1574
rect 16962 1444 16972 1532
rect 17012 1444 17022 1532
rect 16962 1402 17022 1444
rect 17106 1532 17166 1574
rect 17106 1444 17116 1532
rect 17156 1444 17166 1532
rect 17106 1402 17166 1444
rect 17394 1558 17454 1574
rect 17394 1518 17404 1558
rect 17444 1518 17454 1558
rect 17394 1458 17454 1518
rect 17394 1418 17404 1458
rect 17444 1418 17454 1458
rect 17394 1402 17454 1418
rect 17538 1558 17598 1574
rect 17538 1518 17548 1558
rect 17588 1518 17598 1558
rect 17538 1458 17598 1518
rect 17538 1418 17548 1458
rect 17588 1418 17598 1458
rect 17538 1402 17598 1418
rect 17682 1558 17742 1574
rect 17682 1518 17692 1558
rect 17732 1518 17742 1558
rect 17682 1458 17742 1518
rect 17682 1418 17692 1458
rect 17732 1418 17742 1458
rect 17682 1402 17742 1418
rect 17826 1558 17886 1574
rect 17826 1518 17836 1558
rect 17876 1518 17886 1558
rect 17826 1458 17886 1518
rect 17826 1418 17836 1458
rect 17876 1418 17886 1458
rect 17826 1402 17886 1418
rect 17970 1558 18030 1574
rect 17970 1518 17980 1558
rect 18020 1518 18030 1558
rect 17970 1458 18030 1518
rect 17970 1418 17980 1458
rect 18020 1418 18030 1458
rect 17970 1402 18030 1418
rect 18114 1558 18174 1574
rect 18114 1518 18124 1558
rect 18164 1518 18174 1558
rect 18114 1458 18174 1518
rect 18114 1418 18124 1458
rect 18164 1418 18174 1458
rect 18114 1402 18174 1418
rect 18258 1558 18318 1574
rect 18258 1518 18268 1558
rect 18308 1518 18318 1558
rect 18258 1458 18318 1518
rect 18258 1418 18268 1458
rect 18308 1418 18318 1458
rect 18258 1402 18318 1418
rect 18402 1558 18462 1574
rect 18402 1518 18412 1558
rect 18452 1518 18462 1558
rect 18402 1458 18462 1518
rect 18402 1418 18412 1458
rect 18452 1418 18462 1458
rect 18402 1402 18462 1418
rect 18546 1558 18606 1574
rect 18546 1518 18556 1558
rect 18596 1518 18606 1558
rect 18546 1458 18606 1518
rect 18546 1418 18556 1458
rect 18596 1418 18606 1458
rect 18546 1402 18606 1418
rect 18690 1558 18750 1574
rect 18690 1518 18700 1558
rect 18740 1518 18750 1558
rect 18690 1458 18750 1518
rect 18690 1418 18700 1458
rect 18740 1418 18750 1458
rect 18690 1402 18750 1418
rect 18834 1558 18894 1574
rect 18834 1518 18844 1558
rect 18884 1518 18894 1558
rect 18834 1458 18894 1518
rect 18834 1418 18844 1458
rect 18884 1418 18894 1458
rect 18834 1402 18894 1418
rect 18978 1558 19038 1574
rect 18978 1518 18988 1558
rect 19028 1518 19038 1558
rect 18978 1458 19038 1518
rect 18978 1418 18988 1458
rect 19028 1418 19038 1458
rect 18978 1402 19038 1418
rect 19122 1558 19182 1574
rect 19122 1518 19132 1558
rect 19172 1518 19182 1558
rect 19122 1458 19182 1518
rect 19122 1418 19132 1458
rect 19172 1418 19182 1458
rect 19122 1402 19182 1418
rect 19266 1558 19326 1574
rect 19266 1518 19276 1558
rect 19316 1518 19326 1558
rect 19266 1458 19326 1518
rect 19266 1418 19276 1458
rect 19316 1418 19326 1458
rect 19266 1402 19326 1418
rect 19410 1558 19470 1574
rect 19410 1518 19420 1558
rect 19460 1518 19470 1558
rect 19410 1458 19470 1518
rect 19410 1418 19420 1458
rect 19460 1418 19470 1458
rect 19410 1402 19470 1418
rect 19554 1558 19614 1574
rect 19554 1518 19564 1558
rect 19604 1518 19614 1558
rect 19554 1458 19614 1518
rect 19554 1418 19564 1458
rect 19604 1418 19614 1458
rect 19554 1402 19614 1418
rect 19698 1558 19758 1574
rect 19698 1518 19708 1558
rect 19748 1518 19758 1558
rect 19698 1458 19758 1518
rect 19698 1418 19708 1458
rect 19748 1418 19758 1458
rect 19698 1402 19758 1418
rect 19842 1558 19902 1574
rect 19842 1518 19852 1558
rect 19892 1518 19902 1558
rect 19842 1458 19902 1518
rect 19842 1418 19852 1458
rect 19892 1418 19902 1458
rect 19842 1402 19902 1418
rect 19986 1558 20046 1574
rect 19986 1518 19996 1558
rect 20036 1518 20046 1558
rect 19986 1458 20046 1518
rect 19986 1418 19996 1458
rect 20036 1418 20046 1458
rect 19986 1402 20046 1418
rect 20130 1558 20190 1574
rect 20130 1518 20140 1558
rect 20180 1518 20190 1558
rect 20130 1458 20190 1518
rect 20130 1418 20140 1458
rect 20180 1418 20190 1458
rect 20130 1402 20190 1418
rect 20274 1558 20334 1574
rect 20274 1518 20284 1558
rect 20324 1518 20334 1558
rect 20274 1458 20334 1518
rect 20274 1418 20284 1458
rect 20324 1418 20334 1458
rect 20274 1402 20334 1418
rect 20418 1558 20478 1574
rect 20418 1518 20428 1558
rect 20468 1518 20478 1558
rect 20418 1458 20478 1518
rect 20418 1418 20428 1458
rect 20468 1418 20478 1458
rect 20418 1402 20478 1418
rect 20562 1558 20622 1574
rect 20562 1518 20572 1558
rect 20612 1518 20622 1558
rect 20562 1458 20622 1518
rect 20562 1418 20572 1458
rect 20612 1418 20622 1458
rect 20562 1402 20622 1418
rect 20706 1558 20766 1574
rect 20706 1518 20716 1558
rect 20756 1518 20766 1558
rect 20706 1458 20766 1518
rect 20706 1418 20716 1458
rect 20756 1418 20766 1458
rect 20706 1402 20766 1418
rect 20850 1558 20910 1574
rect 20850 1518 20860 1558
rect 20900 1518 20910 1558
rect 20850 1458 20910 1518
rect 20850 1418 20860 1458
rect 20900 1418 20910 1458
rect 20850 1402 20910 1418
rect 776 1313 950 1332
rect 776 1279 796 1313
rect 830 1279 904 1313
rect 938 1279 950 1313
rect 776 1260 950 1279
rect 1352 1313 1526 1332
rect 1352 1279 1372 1313
rect 1406 1279 1480 1313
rect 1514 1279 1526 1313
rect 1352 1260 1526 1279
rect 1928 1313 2102 1332
rect 1928 1279 1948 1313
rect 1982 1279 2056 1313
rect 2090 1279 2102 1313
rect 1928 1260 2102 1279
rect 3080 1313 3254 1332
rect 3080 1279 3100 1313
rect 3134 1279 3208 1313
rect 3242 1279 3254 1313
rect 3080 1260 3254 1279
rect 3656 1313 3830 1332
rect 3656 1279 3676 1313
rect 3710 1279 3784 1313
rect 3818 1279 3830 1313
rect 3656 1260 3830 1279
rect 4232 1313 4406 1332
rect 4232 1279 4252 1313
rect 4286 1279 4360 1313
rect 4394 1279 4406 1313
rect 4232 1260 4406 1279
rect 5960 1313 6134 1332
rect 5960 1279 5980 1313
rect 6014 1279 6088 1313
rect 6122 1279 6134 1313
rect 5960 1260 6134 1279
rect 6536 1313 6710 1332
rect 6536 1279 6556 1313
rect 6590 1279 6664 1313
rect 6698 1279 6710 1313
rect 6536 1260 6710 1279
rect 7112 1313 7286 1332
rect 7112 1279 7132 1313
rect 7166 1279 7240 1313
rect 7274 1279 7286 1313
rect 7112 1260 7286 1279
rect 7688 1313 7862 1332
rect 7688 1279 7708 1313
rect 7742 1279 7816 1313
rect 7850 1279 7862 1313
rect 7688 1260 7862 1279
rect 8174 1314 8264 1332
rect 8174 1278 8196 1314
rect 8232 1278 8264 1314
rect 8174 1260 8264 1278
rect 8438 1314 8528 1332
rect 8438 1278 8474 1314
rect 8510 1278 8528 1314
rect 8438 1260 8528 1278
rect 9416 1313 9590 1332
rect 9416 1279 9436 1313
rect 9470 1279 9544 1313
rect 9578 1279 9590 1313
rect 9416 1260 9590 1279
rect 9992 1313 10166 1332
rect 9992 1279 10012 1313
rect 10046 1279 10120 1313
rect 10154 1279 10166 1313
rect 9992 1260 10166 1279
rect 10568 1313 10742 1332
rect 10568 1279 10588 1313
rect 10622 1279 10696 1313
rect 10730 1279 10742 1313
rect 10568 1260 10742 1279
rect 11054 1314 11144 1332
rect 11054 1278 11076 1314
rect 11112 1278 11144 1314
rect 11054 1260 11144 1278
rect 11318 1314 11408 1332
rect 11318 1278 11354 1314
rect 11390 1278 11408 1314
rect 11318 1260 11408 1278
rect 12008 1313 12182 1332
rect 12008 1279 12028 1313
rect 12062 1279 12136 1313
rect 12170 1279 12182 1313
rect 12008 1260 12182 1279
rect 12584 1313 12758 1332
rect 12584 1279 12604 1313
rect 12638 1279 12712 1313
rect 12746 1279 12758 1313
rect 12584 1260 12758 1279
rect 13160 1313 13334 1332
rect 13160 1279 13180 1313
rect 13214 1279 13288 1313
rect 13322 1279 13334 1313
rect 13160 1260 13334 1279
rect 13736 1313 13910 1332
rect 13736 1279 13756 1313
rect 13790 1279 13864 1313
rect 13898 1279 13910 1313
rect 13736 1260 13910 1279
rect 14888 1313 15062 1332
rect 14888 1279 14908 1313
rect 14942 1279 15016 1313
rect 15050 1279 15062 1313
rect 14888 1260 15062 1279
rect 15466 1313 15640 1332
rect 15466 1279 15478 1313
rect 15512 1279 15586 1313
rect 15620 1279 15640 1313
rect 15466 1260 15640 1279
rect 16040 1313 16214 1332
rect 16040 1279 16060 1313
rect 16094 1279 16168 1313
rect 16202 1279 16214 1313
rect 16040 1260 16214 1279
rect 16328 1313 16502 1332
rect 16328 1279 16348 1313
rect 16382 1279 16456 1313
rect 16490 1279 16502 1313
rect 16328 1260 16502 1279
rect 17480 1313 17654 1332
rect 17480 1279 17500 1313
rect 17534 1279 17608 1313
rect 17642 1279 17654 1313
rect 17480 1260 17654 1279
rect 17768 1313 17942 1332
rect 17768 1279 17788 1313
rect 17822 1279 17896 1313
rect 17930 1279 17942 1313
rect 17768 1260 17942 1279
rect 18056 1313 18230 1332
rect 18056 1279 18076 1313
rect 18110 1279 18184 1313
rect 18218 1279 18230 1313
rect 18056 1260 18230 1279
rect 18344 1313 18518 1332
rect 18344 1279 18364 1313
rect 18398 1279 18472 1313
rect 18506 1279 18518 1313
rect 18344 1260 18518 1279
rect 18632 1313 18806 1332
rect 18632 1279 18652 1313
rect 18686 1279 18760 1313
rect 18794 1279 18806 1313
rect 18632 1260 18806 1279
rect 18920 1313 19094 1332
rect 18920 1279 18940 1313
rect 18974 1279 19048 1313
rect 19082 1279 19094 1313
rect 18920 1260 19094 1279
rect 19208 1313 19382 1332
rect 19208 1279 19228 1313
rect 19262 1279 19336 1313
rect 19370 1279 19382 1313
rect 19208 1260 19382 1279
rect 19496 1313 19670 1332
rect 19496 1279 19516 1313
rect 19550 1279 19624 1313
rect 19658 1279 19670 1313
rect 19496 1260 19670 1279
rect 19784 1313 19958 1332
rect 19784 1279 19804 1313
rect 19838 1279 19912 1313
rect 19946 1279 19958 1313
rect 19784 1260 19958 1279
rect 20072 1313 20246 1332
rect 20072 1279 20092 1313
rect 20126 1279 20200 1313
rect 20234 1279 20246 1313
rect 20072 1260 20246 1279
rect 20360 1313 20534 1332
rect 20360 1279 20380 1313
rect 20414 1279 20488 1313
rect 20522 1279 20534 1313
rect 20360 1260 20534 1279
rect 20648 1313 20822 1332
rect 20648 1279 20668 1313
rect 20702 1279 20776 1313
rect 20810 1279 20822 1313
rect 20648 1260 20822 1279
rect 776 737 950 756
rect 776 703 796 737
rect 830 703 904 737
rect 938 703 950 737
rect 776 684 950 703
rect 1352 737 1526 756
rect 1352 703 1372 737
rect 1406 703 1480 737
rect 1514 703 1526 737
rect 1352 684 1526 703
rect 1928 737 2102 756
rect 1928 703 1948 737
rect 1982 703 2056 737
rect 2090 703 2102 737
rect 1928 684 2102 703
rect 3080 737 3254 756
rect 3080 703 3100 737
rect 3134 703 3208 737
rect 3242 703 3254 737
rect 3080 684 3254 703
rect 3656 737 3830 756
rect 3656 703 3676 737
rect 3710 703 3784 737
rect 3818 703 3830 737
rect 3656 684 3830 703
rect 4232 737 4406 756
rect 4232 703 4252 737
rect 4286 703 4360 737
rect 4394 703 4406 737
rect 4232 684 4406 703
rect 5960 737 6134 756
rect 5960 703 5980 737
rect 6014 703 6088 737
rect 6122 703 6134 737
rect 5960 684 6134 703
rect 6536 737 6710 756
rect 6536 703 6556 737
rect 6590 703 6664 737
rect 6698 703 6710 737
rect 6536 684 6710 703
rect 7112 737 7286 756
rect 7112 703 7132 737
rect 7166 703 7240 737
rect 7274 703 7286 737
rect 7112 684 7286 703
rect 7688 737 7862 756
rect 7688 703 7708 737
rect 7742 703 7816 737
rect 7850 703 7862 737
rect 7688 684 7862 703
rect 8174 738 8264 756
rect 8174 702 8196 738
rect 8232 702 8264 738
rect 8174 684 8264 702
rect 8438 738 8528 756
rect 8438 702 8480 738
rect 8516 702 8528 738
rect 8438 684 8528 702
rect 9416 737 9590 756
rect 9416 703 9436 737
rect 9470 703 9544 737
rect 9578 703 9590 737
rect 9416 684 9590 703
rect 9992 737 10166 756
rect 9992 703 10012 737
rect 10046 703 10120 737
rect 10154 703 10166 737
rect 9992 684 10166 703
rect 10568 737 10742 756
rect 10568 703 10588 737
rect 10622 703 10696 737
rect 10730 703 10742 737
rect 10568 684 10742 703
rect 11054 738 11144 756
rect 11054 702 11076 738
rect 11112 702 11144 738
rect 11054 684 11144 702
rect 11318 738 11408 756
rect 11318 702 11360 738
rect 11396 702 11408 738
rect 11318 684 11408 702
rect 12008 737 12182 756
rect 12008 703 12028 737
rect 12062 703 12136 737
rect 12170 703 12182 737
rect 12008 684 12182 703
rect 12584 737 12758 756
rect 12584 703 12604 737
rect 12638 703 12712 737
rect 12746 703 12758 737
rect 12584 684 12758 703
rect 13160 737 13334 756
rect 13160 703 13180 737
rect 13214 703 13288 737
rect 13322 703 13334 737
rect 13160 684 13334 703
rect 13736 737 13910 756
rect 13736 703 13756 737
rect 13790 703 13864 737
rect 13898 703 13910 737
rect 13736 684 13910 703
rect 14888 737 15062 756
rect 14888 703 14908 737
rect 14942 703 15016 737
rect 15050 703 15062 737
rect 14888 684 15062 703
rect 15466 737 15640 756
rect 15466 703 15478 737
rect 15512 703 15586 737
rect 15620 703 15640 737
rect 15466 684 15640 703
rect 16040 737 16214 756
rect 16040 703 16060 737
rect 16094 703 16168 737
rect 16202 703 16214 737
rect 16040 684 16214 703
rect 16328 737 16502 756
rect 16328 703 16348 737
rect 16382 703 16456 737
rect 16490 703 16502 737
rect 16328 684 16502 703
rect 17480 737 17654 756
rect 17480 703 17500 737
rect 17534 703 17608 737
rect 17642 703 17654 737
rect 17480 684 17654 703
rect 17768 737 17942 756
rect 17768 703 17788 737
rect 17822 703 17896 737
rect 17930 703 17942 737
rect 17768 684 17942 703
rect 18056 737 18230 756
rect 18056 703 18076 737
rect 18110 703 18184 737
rect 18218 703 18230 737
rect 18056 684 18230 703
rect 18344 737 18518 756
rect 18344 703 18364 737
rect 18398 703 18472 737
rect 18506 703 18518 737
rect 18344 684 18518 703
rect 18632 737 18806 756
rect 18632 703 18652 737
rect 18686 703 18760 737
rect 18794 703 18806 737
rect 18632 684 18806 703
rect 18920 737 19094 756
rect 18920 703 18940 737
rect 18974 703 19048 737
rect 19082 703 19094 737
rect 18920 684 19094 703
rect 19208 737 19382 756
rect 19208 703 19228 737
rect 19262 703 19336 737
rect 19370 703 19382 737
rect 19208 684 19382 703
rect 19496 737 19670 756
rect 19496 703 19516 737
rect 19550 703 19624 737
rect 19658 703 19670 737
rect 19496 684 19670 703
rect 19784 737 19958 756
rect 19784 703 19804 737
rect 19838 703 19912 737
rect 19946 703 19958 737
rect 19784 684 19958 703
rect 20072 737 20246 756
rect 20072 703 20092 737
rect 20126 703 20200 737
rect 20234 703 20246 737
rect 20072 684 20246 703
rect 20360 737 20534 756
rect 20360 703 20380 737
rect 20414 703 20488 737
rect 20522 703 20534 737
rect 20360 684 20534 703
rect 20648 737 20822 756
rect 20648 703 20668 737
rect 20702 703 20776 737
rect 20810 703 20822 737
rect 20648 684 20822 703
rect 690 578 750 594
rect 690 538 700 578
rect 740 538 750 578
rect 114 480 174 504
rect 114 328 124 480
rect 164 328 174 480
rect 114 304 174 328
rect 258 480 318 504
rect 258 328 268 480
rect 308 328 318 480
rect 258 304 318 328
rect 402 480 462 504
rect 402 328 412 480
rect 452 328 462 480
rect 402 304 462 328
rect 690 478 750 538
rect 690 438 700 478
rect 740 438 750 478
rect 690 378 750 438
rect 690 338 700 378
rect 740 338 750 378
rect 690 278 750 338
rect 690 238 700 278
rect 740 238 750 278
rect 690 222 750 238
rect 834 578 894 594
rect 834 538 844 578
rect 884 538 894 578
rect 834 478 894 538
rect 834 438 844 478
rect 884 438 894 478
rect 834 378 894 438
rect 834 338 844 378
rect 884 338 894 378
rect 834 278 894 338
rect 834 238 844 278
rect 884 238 894 278
rect 834 222 894 238
rect 978 578 1038 594
rect 978 538 988 578
rect 1028 538 1038 578
rect 978 478 1038 538
rect 978 438 988 478
rect 1028 438 1038 478
rect 978 378 1038 438
rect 978 338 988 378
rect 1028 338 1038 378
rect 978 278 1038 338
rect 978 238 988 278
rect 1028 238 1038 278
rect 978 222 1038 238
rect 1266 578 1326 594
rect 1266 538 1276 578
rect 1316 538 1326 578
rect 1266 478 1326 538
rect 1266 438 1276 478
rect 1316 438 1326 478
rect 1266 378 1326 438
rect 1266 338 1276 378
rect 1316 338 1326 378
rect 1266 278 1326 338
rect 1266 238 1276 278
rect 1316 238 1326 278
rect 1266 222 1326 238
rect 1410 578 1470 594
rect 1410 538 1420 578
rect 1460 538 1470 578
rect 1410 478 1470 538
rect 1410 438 1420 478
rect 1460 438 1470 478
rect 1410 378 1470 438
rect 1410 338 1420 378
rect 1460 338 1470 378
rect 1410 278 1470 338
rect 1410 238 1420 278
rect 1460 238 1470 278
rect 1410 222 1470 238
rect 1554 578 1614 594
rect 1554 538 1564 578
rect 1604 538 1614 578
rect 1554 478 1614 538
rect 1554 438 1564 478
rect 1604 438 1614 478
rect 1554 378 1614 438
rect 1554 338 1564 378
rect 1604 338 1614 378
rect 1554 278 1614 338
rect 1554 238 1564 278
rect 1604 238 1614 278
rect 1554 222 1614 238
rect 1842 578 1902 594
rect 1842 538 1852 578
rect 1892 538 1902 578
rect 1842 478 1902 538
rect 1842 438 1852 478
rect 1892 438 1902 478
rect 1842 378 1902 438
rect 1842 338 1852 378
rect 1892 338 1902 378
rect 1842 278 1902 338
rect 1842 238 1852 278
rect 1892 238 1902 278
rect 1842 222 1902 238
rect 1986 578 2046 594
rect 1986 538 1996 578
rect 2036 538 2046 578
rect 1986 478 2046 538
rect 1986 438 1996 478
rect 2036 438 2046 478
rect 1986 378 2046 438
rect 1986 338 1996 378
rect 2036 338 2046 378
rect 1986 278 2046 338
rect 1986 238 1996 278
rect 2036 238 2046 278
rect 1986 222 2046 238
rect 2130 578 2190 594
rect 2130 538 2140 578
rect 2180 538 2190 578
rect 2130 478 2190 538
rect 2130 438 2140 478
rect 2180 438 2190 478
rect 2130 378 2190 438
rect 2130 338 2140 378
rect 2180 338 2190 378
rect 2130 278 2190 338
rect 2130 238 2140 278
rect 2180 238 2190 278
rect 2130 222 2190 238
rect 2994 578 3054 594
rect 2994 538 3004 578
rect 3044 538 3054 578
rect 2994 478 3054 538
rect 2994 438 3004 478
rect 3044 438 3054 478
rect 2994 378 3054 438
rect 2994 338 3004 378
rect 3044 338 3054 378
rect 2994 278 3054 338
rect 2994 238 3004 278
rect 3044 238 3054 278
rect 2994 222 3054 238
rect 3138 578 3198 594
rect 3138 538 3148 578
rect 3188 538 3198 578
rect 3138 478 3198 538
rect 3138 438 3148 478
rect 3188 438 3198 478
rect 3138 378 3198 438
rect 3138 338 3148 378
rect 3188 338 3198 378
rect 3138 278 3198 338
rect 3138 238 3148 278
rect 3188 238 3198 278
rect 3138 222 3198 238
rect 3282 578 3342 594
rect 3282 538 3292 578
rect 3332 538 3342 578
rect 3282 478 3342 538
rect 3282 438 3292 478
rect 3332 438 3342 478
rect 3282 378 3342 438
rect 3282 338 3292 378
rect 3332 338 3342 378
rect 3282 278 3342 338
rect 3282 238 3292 278
rect 3332 238 3342 278
rect 3282 222 3342 238
rect 3570 578 3630 594
rect 3570 538 3580 578
rect 3620 538 3630 578
rect 3570 478 3630 538
rect 3570 438 3580 478
rect 3620 438 3630 478
rect 3570 378 3630 438
rect 3570 338 3580 378
rect 3620 338 3630 378
rect 3570 278 3630 338
rect 3570 238 3580 278
rect 3620 238 3630 278
rect 3570 222 3630 238
rect 3714 578 3774 594
rect 3714 538 3724 578
rect 3764 538 3774 578
rect 3714 478 3774 538
rect 3714 438 3724 478
rect 3764 438 3774 478
rect 3714 378 3774 438
rect 3714 338 3724 378
rect 3764 338 3774 378
rect 3714 278 3774 338
rect 3714 238 3724 278
rect 3764 238 3774 278
rect 3714 222 3774 238
rect 3858 578 3918 594
rect 3858 538 3868 578
rect 3908 538 3918 578
rect 3858 478 3918 538
rect 3858 438 3868 478
rect 3908 438 3918 478
rect 3858 378 3918 438
rect 3858 338 3868 378
rect 3908 338 3918 378
rect 3858 278 3918 338
rect 3858 238 3868 278
rect 3908 238 3918 278
rect 3858 222 3918 238
rect 4146 578 4206 594
rect 4146 538 4156 578
rect 4196 538 4206 578
rect 4146 478 4206 538
rect 4146 438 4156 478
rect 4196 438 4206 478
rect 4146 378 4206 438
rect 4146 338 4156 378
rect 4196 338 4206 378
rect 4146 278 4206 338
rect 4146 238 4156 278
rect 4196 238 4206 278
rect 4146 222 4206 238
rect 4290 578 4350 594
rect 4290 538 4300 578
rect 4340 538 4350 578
rect 4290 478 4350 538
rect 4290 438 4300 478
rect 4340 438 4350 478
rect 4290 378 4350 438
rect 4290 338 4300 378
rect 4340 338 4350 378
rect 4290 278 4350 338
rect 4290 238 4300 278
rect 4340 238 4350 278
rect 4290 222 4350 238
rect 4434 578 4494 594
rect 4434 538 4444 578
rect 4484 538 4494 578
rect 4434 478 4494 538
rect 5874 578 5934 594
rect 5874 538 5884 578
rect 5924 538 5934 578
rect 4434 438 4444 478
rect 4484 438 4494 478
rect 4434 378 4494 438
rect 4434 338 4444 378
rect 4484 338 4494 378
rect 4434 278 4494 338
rect 4722 480 4782 504
rect 4722 328 4732 480
rect 4772 328 4782 480
rect 4722 304 4782 328
rect 4866 480 4926 504
rect 4866 328 4876 480
rect 4916 328 4926 480
rect 4866 304 4926 328
rect 5010 480 5070 504
rect 5010 328 5020 480
rect 5060 328 5070 480
rect 5010 304 5070 328
rect 5298 480 5358 504
rect 5298 328 5308 480
rect 5348 328 5358 480
rect 5298 304 5358 328
rect 5442 480 5502 504
rect 5442 328 5452 480
rect 5492 328 5502 480
rect 5442 304 5502 328
rect 5586 480 5646 504
rect 5586 328 5596 480
rect 5636 328 5646 480
rect 5586 304 5646 328
rect 5874 478 5934 538
rect 5874 438 5884 478
rect 5924 438 5934 478
rect 5874 378 5934 438
rect 5874 338 5884 378
rect 5924 338 5934 378
rect 4434 238 4444 278
rect 4484 238 4494 278
rect 4434 222 4494 238
rect 5874 278 5934 338
rect 5874 238 5884 278
rect 5924 238 5934 278
rect 5874 222 5934 238
rect 6018 578 6078 594
rect 6018 538 6028 578
rect 6068 538 6078 578
rect 6018 478 6078 538
rect 6018 438 6028 478
rect 6068 438 6078 478
rect 6018 378 6078 438
rect 6018 338 6028 378
rect 6068 338 6078 378
rect 6018 278 6078 338
rect 6018 238 6028 278
rect 6068 238 6078 278
rect 6018 222 6078 238
rect 6162 578 6222 594
rect 6162 538 6172 578
rect 6212 538 6222 578
rect 6162 478 6222 538
rect 6162 438 6172 478
rect 6212 438 6222 478
rect 6162 378 6222 438
rect 6162 338 6172 378
rect 6212 338 6222 378
rect 6162 278 6222 338
rect 6162 238 6172 278
rect 6212 238 6222 278
rect 6162 222 6222 238
rect 6450 578 6510 594
rect 6450 538 6460 578
rect 6500 538 6510 578
rect 6450 478 6510 538
rect 6450 438 6460 478
rect 6500 438 6510 478
rect 6450 378 6510 438
rect 6450 338 6460 378
rect 6500 338 6510 378
rect 6450 278 6510 338
rect 6450 238 6460 278
rect 6500 238 6510 278
rect 6450 222 6510 238
rect 6594 578 6654 594
rect 6594 538 6604 578
rect 6644 538 6654 578
rect 6594 478 6654 538
rect 6594 438 6604 478
rect 6644 438 6654 478
rect 6594 378 6654 438
rect 6594 338 6604 378
rect 6644 338 6654 378
rect 6594 278 6654 338
rect 6594 238 6604 278
rect 6644 238 6654 278
rect 6594 222 6654 238
rect 6738 578 6798 594
rect 6738 538 6748 578
rect 6788 538 6798 578
rect 6738 478 6798 538
rect 6738 438 6748 478
rect 6788 438 6798 478
rect 6738 378 6798 438
rect 6738 338 6748 378
rect 6788 338 6798 378
rect 6738 278 6798 338
rect 6738 238 6748 278
rect 6788 238 6798 278
rect 6738 222 6798 238
rect 7026 578 7086 594
rect 7026 538 7036 578
rect 7076 538 7086 578
rect 7026 478 7086 538
rect 7026 438 7036 478
rect 7076 438 7086 478
rect 7026 378 7086 438
rect 7026 338 7036 378
rect 7076 338 7086 378
rect 7026 278 7086 338
rect 7026 238 7036 278
rect 7076 238 7086 278
rect 7026 222 7086 238
rect 7170 578 7230 594
rect 7170 538 7180 578
rect 7220 538 7230 578
rect 7170 478 7230 538
rect 7170 438 7180 478
rect 7220 438 7230 478
rect 7170 378 7230 438
rect 7170 338 7180 378
rect 7220 338 7230 378
rect 7170 278 7230 338
rect 7170 238 7180 278
rect 7220 238 7230 278
rect 7170 222 7230 238
rect 7314 578 7374 594
rect 7314 538 7324 578
rect 7364 538 7374 578
rect 7314 478 7374 538
rect 7314 438 7324 478
rect 7364 438 7374 478
rect 7314 378 7374 438
rect 7314 338 7324 378
rect 7364 338 7374 378
rect 7314 278 7374 338
rect 7314 238 7324 278
rect 7364 238 7374 278
rect 7314 222 7374 238
rect 7602 578 7662 594
rect 7602 538 7612 578
rect 7652 538 7662 578
rect 7602 478 7662 538
rect 7602 438 7612 478
rect 7652 438 7662 478
rect 7602 378 7662 438
rect 7602 338 7612 378
rect 7652 338 7662 378
rect 7602 278 7662 338
rect 7602 238 7612 278
rect 7652 238 7662 278
rect 7602 222 7662 238
rect 7746 578 7806 594
rect 7746 538 7756 578
rect 7796 538 7806 578
rect 7746 478 7806 538
rect 7746 438 7756 478
rect 7796 438 7806 478
rect 7746 378 7806 438
rect 7746 338 7756 378
rect 7796 338 7806 378
rect 7746 278 7806 338
rect 7746 238 7756 278
rect 7796 238 7806 278
rect 7746 222 7806 238
rect 7890 578 7950 594
rect 7890 538 7900 578
rect 7940 538 7950 578
rect 7890 478 7950 538
rect 7890 438 7900 478
rect 7940 438 7950 478
rect 7890 378 7950 438
rect 7890 338 7900 378
rect 7940 338 7950 378
rect 7890 278 7950 338
rect 7890 238 7900 278
rect 7940 238 7950 278
rect 7890 222 7950 238
rect 8178 578 8238 594
rect 8178 538 8188 578
rect 8228 538 8238 578
rect 8178 478 8238 538
rect 8178 438 8188 478
rect 8228 438 8238 478
rect 8178 378 8238 438
rect 8178 338 8188 378
rect 8228 338 8238 378
rect 8178 278 8238 338
rect 8178 238 8188 278
rect 8228 238 8238 278
rect 8178 222 8238 238
rect 8322 578 8382 594
rect 8322 538 8332 578
rect 8372 538 8382 578
rect 8322 478 8382 538
rect 8322 438 8332 478
rect 8372 438 8382 478
rect 8322 378 8382 438
rect 8322 338 8332 378
rect 8372 338 8382 378
rect 8322 278 8382 338
rect 8322 238 8332 278
rect 8372 238 8382 278
rect 8322 222 8382 238
rect 8466 578 8526 594
rect 8466 538 8476 578
rect 8516 538 8526 578
rect 8466 478 8526 538
rect 9330 578 9390 594
rect 9330 538 9340 578
rect 9380 538 9390 578
rect 8466 438 8476 478
rect 8516 438 8526 478
rect 8466 378 8526 438
rect 8466 338 8476 378
rect 8516 338 8526 378
rect 8466 278 8526 338
rect 8754 480 8814 504
rect 8754 328 8764 480
rect 8804 328 8814 480
rect 8754 304 8814 328
rect 8898 480 8958 504
rect 8898 328 8908 480
rect 8948 328 8958 480
rect 8898 304 8958 328
rect 9042 480 9102 504
rect 9042 328 9052 480
rect 9092 328 9102 480
rect 9042 304 9102 328
rect 9330 478 9390 538
rect 9330 438 9340 478
rect 9380 438 9390 478
rect 9330 378 9390 438
rect 9330 338 9340 378
rect 9380 338 9390 378
rect 8466 238 8476 278
rect 8516 238 8526 278
rect 8466 222 8526 238
rect 9330 278 9390 338
rect 9330 238 9340 278
rect 9380 238 9390 278
rect 9330 222 9390 238
rect 9474 578 9534 594
rect 9474 538 9484 578
rect 9524 538 9534 578
rect 9474 478 9534 538
rect 9474 438 9484 478
rect 9524 438 9534 478
rect 9474 378 9534 438
rect 9474 338 9484 378
rect 9524 338 9534 378
rect 9474 278 9534 338
rect 9474 238 9484 278
rect 9524 238 9534 278
rect 9474 222 9534 238
rect 9618 578 9678 594
rect 9618 538 9628 578
rect 9668 538 9678 578
rect 9618 478 9678 538
rect 9618 438 9628 478
rect 9668 438 9678 478
rect 9618 378 9678 438
rect 9618 338 9628 378
rect 9668 338 9678 378
rect 9618 278 9678 338
rect 9618 238 9628 278
rect 9668 238 9678 278
rect 9618 222 9678 238
rect 9906 578 9966 594
rect 9906 538 9916 578
rect 9956 538 9966 578
rect 9906 478 9966 538
rect 9906 438 9916 478
rect 9956 438 9966 478
rect 9906 378 9966 438
rect 9906 338 9916 378
rect 9956 338 9966 378
rect 9906 278 9966 338
rect 9906 238 9916 278
rect 9956 238 9966 278
rect 9906 222 9966 238
rect 10050 578 10110 594
rect 10050 538 10060 578
rect 10100 538 10110 578
rect 10050 478 10110 538
rect 10050 438 10060 478
rect 10100 438 10110 478
rect 10050 378 10110 438
rect 10050 338 10060 378
rect 10100 338 10110 378
rect 10050 278 10110 338
rect 10050 238 10060 278
rect 10100 238 10110 278
rect 10050 222 10110 238
rect 10194 578 10254 594
rect 10194 538 10204 578
rect 10244 538 10254 578
rect 10194 478 10254 538
rect 10194 438 10204 478
rect 10244 438 10254 478
rect 10194 378 10254 438
rect 10194 338 10204 378
rect 10244 338 10254 378
rect 10194 278 10254 338
rect 10194 238 10204 278
rect 10244 238 10254 278
rect 10194 222 10254 238
rect 10482 578 10542 594
rect 10482 538 10492 578
rect 10532 538 10542 578
rect 10482 478 10542 538
rect 10482 438 10492 478
rect 10532 438 10542 478
rect 10482 378 10542 438
rect 10482 338 10492 378
rect 10532 338 10542 378
rect 10482 278 10542 338
rect 10482 238 10492 278
rect 10532 238 10542 278
rect 10482 222 10542 238
rect 10626 578 10686 594
rect 10626 538 10636 578
rect 10676 538 10686 578
rect 10626 478 10686 538
rect 10626 438 10636 478
rect 10676 438 10686 478
rect 10626 378 10686 438
rect 10626 338 10636 378
rect 10676 338 10686 378
rect 10626 278 10686 338
rect 10626 238 10636 278
rect 10676 238 10686 278
rect 10626 222 10686 238
rect 10770 578 10830 594
rect 10770 538 10780 578
rect 10820 538 10830 578
rect 10770 478 10830 538
rect 10770 438 10780 478
rect 10820 438 10830 478
rect 10770 378 10830 438
rect 10770 338 10780 378
rect 10820 338 10830 378
rect 10770 278 10830 338
rect 10770 238 10780 278
rect 10820 238 10830 278
rect 10770 222 10830 238
rect 11058 578 11118 594
rect 11058 538 11068 578
rect 11108 538 11118 578
rect 11058 478 11118 538
rect 11058 438 11068 478
rect 11108 438 11118 478
rect 11058 378 11118 438
rect 11058 338 11068 378
rect 11108 338 11118 378
rect 11058 278 11118 338
rect 11058 238 11068 278
rect 11108 238 11118 278
rect 11058 222 11118 238
rect 11202 578 11262 594
rect 11202 538 11212 578
rect 11252 538 11262 578
rect 11202 478 11262 538
rect 11202 438 11212 478
rect 11252 438 11262 478
rect 11202 378 11262 438
rect 11202 338 11212 378
rect 11252 338 11262 378
rect 11202 278 11262 338
rect 11202 238 11212 278
rect 11252 238 11262 278
rect 11202 222 11262 238
rect 11346 578 11406 594
rect 11346 538 11356 578
rect 11396 538 11406 578
rect 11346 478 11406 538
rect 11346 438 11356 478
rect 11396 438 11406 478
rect 11346 378 11406 438
rect 11346 338 11356 378
rect 11396 338 11406 378
rect 11346 278 11406 338
rect 11346 238 11356 278
rect 11396 238 11406 278
rect 11346 222 11406 238
rect 11922 578 11982 594
rect 11922 538 11932 578
rect 11972 538 11982 578
rect 11922 478 11982 538
rect 11922 438 11932 478
rect 11972 438 11982 478
rect 11922 378 11982 438
rect 11922 338 11932 378
rect 11972 338 11982 378
rect 11922 278 11982 338
rect 11922 238 11932 278
rect 11972 238 11982 278
rect 11922 222 11982 238
rect 12066 578 12126 594
rect 12066 538 12076 578
rect 12116 538 12126 578
rect 12066 478 12126 538
rect 12066 438 12076 478
rect 12116 438 12126 478
rect 12066 378 12126 438
rect 12066 338 12076 378
rect 12116 338 12126 378
rect 12066 278 12126 338
rect 12066 238 12076 278
rect 12116 238 12126 278
rect 12066 222 12126 238
rect 12210 578 12270 594
rect 12210 538 12220 578
rect 12260 538 12270 578
rect 12210 478 12270 538
rect 12210 438 12220 478
rect 12260 438 12270 478
rect 12210 378 12270 438
rect 12210 338 12220 378
rect 12260 338 12270 378
rect 12210 278 12270 338
rect 12210 238 12220 278
rect 12260 238 12270 278
rect 12210 222 12270 238
rect 12498 578 12558 594
rect 12498 538 12508 578
rect 12548 538 12558 578
rect 12498 478 12558 538
rect 12498 438 12508 478
rect 12548 438 12558 478
rect 12498 378 12558 438
rect 12498 338 12508 378
rect 12548 338 12558 378
rect 12498 278 12558 338
rect 12498 238 12508 278
rect 12548 238 12558 278
rect 12498 222 12558 238
rect 12642 578 12702 594
rect 12642 538 12652 578
rect 12692 538 12702 578
rect 12642 478 12702 538
rect 12642 438 12652 478
rect 12692 438 12702 478
rect 12642 378 12702 438
rect 12642 338 12652 378
rect 12692 338 12702 378
rect 12642 278 12702 338
rect 12642 238 12652 278
rect 12692 238 12702 278
rect 12642 222 12702 238
rect 12786 578 12846 594
rect 12786 538 12796 578
rect 12836 538 12846 578
rect 12786 478 12846 538
rect 12786 438 12796 478
rect 12836 438 12846 478
rect 12786 378 12846 438
rect 12786 338 12796 378
rect 12836 338 12846 378
rect 12786 278 12846 338
rect 12786 238 12796 278
rect 12836 238 12846 278
rect 12786 222 12846 238
rect 13074 578 13134 594
rect 13074 538 13084 578
rect 13124 538 13134 578
rect 13074 478 13134 538
rect 13074 438 13084 478
rect 13124 438 13134 478
rect 13074 378 13134 438
rect 13074 338 13084 378
rect 13124 338 13134 378
rect 13074 278 13134 338
rect 13074 238 13084 278
rect 13124 238 13134 278
rect 13074 222 13134 238
rect 13218 578 13278 594
rect 13218 538 13228 578
rect 13268 538 13278 578
rect 13218 478 13278 538
rect 13218 438 13228 478
rect 13268 438 13278 478
rect 13218 378 13278 438
rect 13218 338 13228 378
rect 13268 338 13278 378
rect 13218 278 13278 338
rect 13218 238 13228 278
rect 13268 238 13278 278
rect 13218 222 13278 238
rect 13362 578 13422 594
rect 13362 538 13372 578
rect 13412 538 13422 578
rect 13362 478 13422 538
rect 13362 438 13372 478
rect 13412 438 13422 478
rect 13362 378 13422 438
rect 13362 338 13372 378
rect 13412 338 13422 378
rect 13362 278 13422 338
rect 13362 238 13372 278
rect 13412 238 13422 278
rect 13362 222 13422 238
rect 13650 578 13710 594
rect 13650 538 13660 578
rect 13700 538 13710 578
rect 13650 478 13710 538
rect 13650 438 13660 478
rect 13700 438 13710 478
rect 13650 378 13710 438
rect 13650 338 13660 378
rect 13700 338 13710 378
rect 13650 278 13710 338
rect 13650 238 13660 278
rect 13700 238 13710 278
rect 13650 222 13710 238
rect 13794 578 13854 594
rect 13794 538 13804 578
rect 13844 538 13854 578
rect 13794 478 13854 538
rect 13794 438 13804 478
rect 13844 438 13854 478
rect 13794 378 13854 438
rect 13794 338 13804 378
rect 13844 338 13854 378
rect 13794 278 13854 338
rect 13794 238 13804 278
rect 13844 238 13854 278
rect 13794 222 13854 238
rect 13938 578 13998 594
rect 13938 538 13948 578
rect 13988 538 13998 578
rect 13938 478 13998 538
rect 14802 578 14862 594
rect 14802 538 14812 578
rect 14852 538 14862 578
rect 13938 438 13948 478
rect 13988 438 13998 478
rect 13938 378 13998 438
rect 13938 338 13948 378
rect 13988 338 13998 378
rect 13938 278 13998 338
rect 14226 480 14286 504
rect 14226 328 14236 480
rect 14276 328 14286 480
rect 14226 304 14286 328
rect 14370 480 14430 504
rect 14370 328 14380 480
rect 14420 328 14430 480
rect 14370 304 14430 328
rect 14514 480 14574 504
rect 14514 328 14524 480
rect 14564 328 14574 480
rect 14514 304 14574 328
rect 14802 478 14862 538
rect 14802 438 14812 478
rect 14852 438 14862 478
rect 14802 378 14862 438
rect 14802 338 14812 378
rect 14852 338 14862 378
rect 13938 238 13948 278
rect 13988 238 13998 278
rect 13938 222 13998 238
rect 14802 278 14862 338
rect 14802 238 14812 278
rect 14852 238 14862 278
rect 14802 222 14862 238
rect 14946 578 15006 594
rect 14946 538 14956 578
rect 14996 538 15006 578
rect 14946 478 15006 538
rect 14946 438 14956 478
rect 14996 438 15006 478
rect 14946 378 15006 438
rect 14946 338 14956 378
rect 14996 338 15006 378
rect 14946 278 15006 338
rect 14946 238 14956 278
rect 14996 238 15006 278
rect 14946 222 15006 238
rect 15090 578 15150 594
rect 15090 538 15100 578
rect 15140 538 15150 578
rect 15090 478 15150 538
rect 15090 438 15100 478
rect 15140 438 15150 478
rect 15090 378 15150 438
rect 15090 338 15100 378
rect 15140 338 15150 378
rect 15090 278 15150 338
rect 15090 238 15100 278
rect 15140 238 15150 278
rect 15090 222 15150 238
rect 15378 578 15438 594
rect 15378 538 15388 578
rect 15428 538 15438 578
rect 15378 478 15438 538
rect 15378 438 15388 478
rect 15428 438 15438 478
rect 15378 378 15438 438
rect 15378 338 15388 378
rect 15428 338 15438 378
rect 15378 278 15438 338
rect 15378 238 15388 278
rect 15428 238 15438 278
rect 15378 222 15438 238
rect 15522 578 15582 594
rect 15522 538 15532 578
rect 15572 538 15582 578
rect 15522 478 15582 538
rect 15522 438 15532 478
rect 15572 438 15582 478
rect 15522 378 15582 438
rect 15522 338 15532 378
rect 15572 338 15582 378
rect 15522 278 15582 338
rect 15522 238 15532 278
rect 15572 238 15582 278
rect 15522 222 15582 238
rect 15666 578 15726 594
rect 15666 538 15676 578
rect 15716 538 15726 578
rect 15666 478 15726 538
rect 15666 438 15676 478
rect 15716 438 15726 478
rect 15666 378 15726 438
rect 15666 338 15676 378
rect 15716 338 15726 378
rect 15666 278 15726 338
rect 15666 238 15676 278
rect 15716 238 15726 278
rect 15666 222 15726 238
rect 15954 578 16014 594
rect 15954 538 15964 578
rect 16004 538 16014 578
rect 15954 478 16014 538
rect 15954 438 15964 478
rect 16004 438 16014 478
rect 15954 378 16014 438
rect 15954 338 15964 378
rect 16004 338 16014 378
rect 15954 278 16014 338
rect 15954 238 15964 278
rect 16004 238 16014 278
rect 15954 222 16014 238
rect 16098 578 16158 594
rect 16098 538 16108 578
rect 16148 538 16158 578
rect 16098 478 16158 538
rect 16098 438 16108 478
rect 16148 438 16158 478
rect 16098 378 16158 438
rect 16098 338 16108 378
rect 16148 338 16158 378
rect 16098 278 16158 338
rect 16098 238 16108 278
rect 16148 238 16158 278
rect 16098 222 16158 238
rect 16242 578 16302 594
rect 16242 538 16252 578
rect 16292 538 16302 578
rect 16242 478 16302 538
rect 16242 438 16252 478
rect 16292 438 16302 478
rect 16242 378 16302 438
rect 16242 338 16252 378
rect 16292 338 16302 378
rect 16242 278 16302 338
rect 16242 238 16252 278
rect 16292 238 16302 278
rect 16242 222 16302 238
rect 16386 578 16446 594
rect 16386 538 16396 578
rect 16436 538 16446 578
rect 16386 478 16446 538
rect 16386 438 16396 478
rect 16436 438 16446 478
rect 16386 378 16446 438
rect 16386 338 16396 378
rect 16436 338 16446 378
rect 16386 278 16446 338
rect 16386 238 16396 278
rect 16436 238 16446 278
rect 16386 222 16446 238
rect 16530 578 16590 594
rect 16530 538 16540 578
rect 16580 538 16590 578
rect 16530 478 16590 538
rect 17394 578 17454 594
rect 17394 538 17404 578
rect 17444 538 17454 578
rect 16530 438 16540 478
rect 16580 438 16590 478
rect 16530 378 16590 438
rect 16530 338 16540 378
rect 16580 338 16590 378
rect 16530 278 16590 338
rect 16818 480 16878 504
rect 16818 328 16828 480
rect 16868 328 16878 480
rect 16818 304 16878 328
rect 16962 480 17022 504
rect 16962 328 16972 480
rect 17012 328 17022 480
rect 16962 304 17022 328
rect 17106 480 17166 504
rect 17106 328 17116 480
rect 17156 328 17166 480
rect 17106 304 17166 328
rect 17394 478 17454 538
rect 17394 438 17404 478
rect 17444 438 17454 478
rect 17394 378 17454 438
rect 17394 338 17404 378
rect 17444 338 17454 378
rect 16530 238 16540 278
rect 16580 238 16590 278
rect 16530 222 16590 238
rect 17394 278 17454 338
rect 17394 238 17404 278
rect 17444 238 17454 278
rect 17394 222 17454 238
rect 17538 578 17598 594
rect 17538 538 17548 578
rect 17588 538 17598 578
rect 17538 478 17598 538
rect 17538 438 17548 478
rect 17588 438 17598 478
rect 17538 378 17598 438
rect 17538 338 17548 378
rect 17588 338 17598 378
rect 17538 278 17598 338
rect 17538 238 17548 278
rect 17588 238 17598 278
rect 17538 222 17598 238
rect 17682 578 17742 594
rect 17682 538 17692 578
rect 17732 538 17742 578
rect 17682 478 17742 538
rect 17682 438 17692 478
rect 17732 438 17742 478
rect 17682 378 17742 438
rect 17682 338 17692 378
rect 17732 338 17742 378
rect 17682 278 17742 338
rect 17682 238 17692 278
rect 17732 238 17742 278
rect 17682 222 17742 238
rect 17826 578 17886 594
rect 17826 538 17836 578
rect 17876 538 17886 578
rect 17826 478 17886 538
rect 17826 438 17836 478
rect 17876 438 17886 478
rect 17826 378 17886 438
rect 17826 338 17836 378
rect 17876 338 17886 378
rect 17826 278 17886 338
rect 17826 238 17836 278
rect 17876 238 17886 278
rect 17826 222 17886 238
rect 17970 578 18030 594
rect 17970 538 17980 578
rect 18020 538 18030 578
rect 17970 478 18030 538
rect 17970 438 17980 478
rect 18020 438 18030 478
rect 17970 378 18030 438
rect 17970 338 17980 378
rect 18020 338 18030 378
rect 17970 278 18030 338
rect 17970 238 17980 278
rect 18020 238 18030 278
rect 17970 222 18030 238
rect 18114 578 18174 594
rect 18114 538 18124 578
rect 18164 538 18174 578
rect 18114 478 18174 538
rect 18114 438 18124 478
rect 18164 438 18174 478
rect 18114 378 18174 438
rect 18114 338 18124 378
rect 18164 338 18174 378
rect 18114 278 18174 338
rect 18114 238 18124 278
rect 18164 238 18174 278
rect 18114 222 18174 238
rect 18258 578 18318 594
rect 18258 538 18268 578
rect 18308 538 18318 578
rect 18258 478 18318 538
rect 18258 438 18268 478
rect 18308 438 18318 478
rect 18258 378 18318 438
rect 18258 338 18268 378
rect 18308 338 18318 378
rect 18258 278 18318 338
rect 18258 238 18268 278
rect 18308 238 18318 278
rect 18258 222 18318 238
rect 18402 578 18462 594
rect 18402 538 18412 578
rect 18452 538 18462 578
rect 18402 478 18462 538
rect 18402 438 18412 478
rect 18452 438 18462 478
rect 18402 378 18462 438
rect 18402 338 18412 378
rect 18452 338 18462 378
rect 18402 278 18462 338
rect 18402 238 18412 278
rect 18452 238 18462 278
rect 18402 222 18462 238
rect 18546 578 18606 594
rect 18546 538 18556 578
rect 18596 538 18606 578
rect 18546 478 18606 538
rect 18546 438 18556 478
rect 18596 438 18606 478
rect 18546 378 18606 438
rect 18546 338 18556 378
rect 18596 338 18606 378
rect 18546 278 18606 338
rect 18546 238 18556 278
rect 18596 238 18606 278
rect 18546 222 18606 238
rect 18690 578 18750 594
rect 18690 538 18700 578
rect 18740 538 18750 578
rect 18690 478 18750 538
rect 18690 438 18700 478
rect 18740 438 18750 478
rect 18690 378 18750 438
rect 18690 338 18700 378
rect 18740 338 18750 378
rect 18690 278 18750 338
rect 18690 238 18700 278
rect 18740 238 18750 278
rect 18690 222 18750 238
rect 18834 578 18894 594
rect 18834 538 18844 578
rect 18884 538 18894 578
rect 18834 478 18894 538
rect 18834 438 18844 478
rect 18884 438 18894 478
rect 18834 378 18894 438
rect 18834 338 18844 378
rect 18884 338 18894 378
rect 18834 278 18894 338
rect 18834 238 18844 278
rect 18884 238 18894 278
rect 18834 222 18894 238
rect 18978 578 19038 594
rect 18978 538 18988 578
rect 19028 538 19038 578
rect 18978 478 19038 538
rect 18978 438 18988 478
rect 19028 438 19038 478
rect 18978 378 19038 438
rect 18978 338 18988 378
rect 19028 338 19038 378
rect 18978 278 19038 338
rect 18978 238 18988 278
rect 19028 238 19038 278
rect 18978 222 19038 238
rect 19122 578 19182 594
rect 19122 538 19132 578
rect 19172 538 19182 578
rect 19122 478 19182 538
rect 19122 438 19132 478
rect 19172 438 19182 478
rect 19122 378 19182 438
rect 19122 338 19132 378
rect 19172 338 19182 378
rect 19122 278 19182 338
rect 19122 238 19132 278
rect 19172 238 19182 278
rect 19122 222 19182 238
rect 19266 578 19326 594
rect 19266 538 19276 578
rect 19316 538 19326 578
rect 19266 478 19326 538
rect 19266 438 19276 478
rect 19316 438 19326 478
rect 19266 378 19326 438
rect 19266 338 19276 378
rect 19316 338 19326 378
rect 19266 278 19326 338
rect 19266 238 19276 278
rect 19316 238 19326 278
rect 19266 222 19326 238
rect 19410 578 19470 594
rect 19410 538 19420 578
rect 19460 538 19470 578
rect 19410 478 19470 538
rect 19410 438 19420 478
rect 19460 438 19470 478
rect 19410 378 19470 438
rect 19410 338 19420 378
rect 19460 338 19470 378
rect 19410 278 19470 338
rect 19410 238 19420 278
rect 19460 238 19470 278
rect 19410 222 19470 238
rect 19554 578 19614 594
rect 19554 538 19564 578
rect 19604 538 19614 578
rect 19554 478 19614 538
rect 19554 438 19564 478
rect 19604 438 19614 478
rect 19554 378 19614 438
rect 19554 338 19564 378
rect 19604 338 19614 378
rect 19554 278 19614 338
rect 19554 238 19564 278
rect 19604 238 19614 278
rect 19554 222 19614 238
rect 19698 578 19758 594
rect 19698 538 19708 578
rect 19748 538 19758 578
rect 19698 478 19758 538
rect 19698 438 19708 478
rect 19748 438 19758 478
rect 19698 378 19758 438
rect 19698 338 19708 378
rect 19748 338 19758 378
rect 19698 278 19758 338
rect 19698 238 19708 278
rect 19748 238 19758 278
rect 19698 222 19758 238
rect 19842 578 19902 594
rect 19842 538 19852 578
rect 19892 538 19902 578
rect 19842 478 19902 538
rect 19842 438 19852 478
rect 19892 438 19902 478
rect 19842 378 19902 438
rect 19842 338 19852 378
rect 19892 338 19902 378
rect 19842 278 19902 338
rect 19842 238 19852 278
rect 19892 238 19902 278
rect 19842 222 19902 238
rect 19986 578 20046 594
rect 19986 538 19996 578
rect 20036 538 20046 578
rect 19986 478 20046 538
rect 19986 438 19996 478
rect 20036 438 20046 478
rect 19986 378 20046 438
rect 19986 338 19996 378
rect 20036 338 20046 378
rect 19986 278 20046 338
rect 19986 238 19996 278
rect 20036 238 20046 278
rect 19986 222 20046 238
rect 20130 578 20190 594
rect 20130 538 20140 578
rect 20180 538 20190 578
rect 20130 478 20190 538
rect 20130 438 20140 478
rect 20180 438 20190 478
rect 20130 378 20190 438
rect 20130 338 20140 378
rect 20180 338 20190 378
rect 20130 278 20190 338
rect 20130 238 20140 278
rect 20180 238 20190 278
rect 20130 222 20190 238
rect 20274 578 20334 594
rect 20274 538 20284 578
rect 20324 538 20334 578
rect 20274 478 20334 538
rect 20274 438 20284 478
rect 20324 438 20334 478
rect 20274 378 20334 438
rect 20274 338 20284 378
rect 20324 338 20334 378
rect 20274 278 20334 338
rect 20274 238 20284 278
rect 20324 238 20334 278
rect 20274 222 20334 238
rect 20418 578 20478 594
rect 20418 538 20428 578
rect 20468 538 20478 578
rect 20418 478 20478 538
rect 20418 438 20428 478
rect 20468 438 20478 478
rect 20418 378 20478 438
rect 20418 338 20428 378
rect 20468 338 20478 378
rect 20418 278 20478 338
rect 20418 238 20428 278
rect 20468 238 20478 278
rect 20418 222 20478 238
rect 20562 578 20622 594
rect 20562 538 20572 578
rect 20612 538 20622 578
rect 20562 478 20622 538
rect 20562 438 20572 478
rect 20612 438 20622 478
rect 20562 378 20622 438
rect 20562 338 20572 378
rect 20612 338 20622 378
rect 20562 278 20622 338
rect 20562 238 20572 278
rect 20612 238 20622 278
rect 20562 222 20622 238
rect 20706 578 20766 594
rect 20706 538 20716 578
rect 20756 538 20766 578
rect 20706 478 20766 538
rect 20706 438 20716 478
rect 20756 438 20766 478
rect 20706 378 20766 438
rect 20706 338 20716 378
rect 20756 338 20766 378
rect 20706 278 20766 338
rect 20706 238 20716 278
rect 20756 238 20766 278
rect 20706 222 20766 238
rect 20850 578 20910 594
rect 20850 538 20860 578
rect 20900 538 20910 578
rect 20850 478 20910 538
rect 20850 438 20860 478
rect 20900 438 20910 478
rect 20850 378 20910 438
rect 20850 338 20860 378
rect 20900 338 20910 378
rect 20850 278 20910 338
rect 20850 238 20860 278
rect 20900 238 20910 278
rect 20850 222 20910 238
<< viali >>
rect 700 3754 740 3794
rect 124 3552 164 3704
rect 268 3552 308 3704
rect 412 3552 452 3704
rect 700 3654 740 3694
rect 700 3554 740 3594
rect 700 3454 740 3494
rect 844 3754 884 3794
rect 844 3654 884 3694
rect 844 3554 884 3594
rect 844 3454 884 3494
rect 988 3754 1028 3794
rect 988 3654 1028 3694
rect 988 3554 1028 3594
rect 988 3454 1028 3494
rect 1276 3754 1316 3794
rect 1276 3654 1316 3694
rect 1276 3554 1316 3594
rect 1276 3454 1316 3494
rect 1420 3754 1460 3794
rect 1420 3654 1460 3694
rect 1420 3554 1460 3594
rect 1420 3454 1460 3494
rect 1564 3754 1604 3794
rect 1564 3654 1604 3694
rect 1564 3554 1604 3594
rect 1564 3454 1604 3494
rect 1852 3754 1892 3794
rect 1852 3654 1892 3694
rect 1852 3554 1892 3594
rect 1852 3454 1892 3494
rect 1996 3754 2036 3794
rect 1996 3654 2036 3694
rect 1996 3554 2036 3594
rect 1996 3454 2036 3494
rect 2140 3754 2180 3794
rect 2140 3654 2180 3694
rect 2140 3554 2180 3594
rect 2140 3454 2180 3494
rect 2428 3754 2468 3794
rect 2428 3654 2468 3694
rect 2428 3554 2468 3594
rect 2428 3454 2468 3494
rect 2572 3754 2612 3794
rect 2572 3654 2612 3694
rect 2572 3554 2612 3594
rect 2572 3454 2612 3494
rect 2716 3754 2756 3794
rect 2716 3654 2756 3694
rect 2716 3554 2756 3594
rect 2716 3454 2756 3494
rect 3004 3754 3044 3794
rect 3004 3654 3044 3694
rect 3004 3554 3044 3594
rect 3004 3454 3044 3494
rect 3148 3754 3188 3794
rect 3148 3654 3188 3694
rect 3148 3554 3188 3594
rect 3148 3454 3188 3494
rect 3292 3754 3332 3794
rect 4156 3754 4196 3794
rect 3292 3654 3332 3694
rect 3292 3554 3332 3594
rect 3580 3552 3620 3704
rect 3724 3552 3764 3704
rect 3868 3552 3908 3704
rect 4156 3654 4196 3694
rect 4156 3554 4196 3594
rect 3292 3454 3332 3494
rect 4156 3454 4196 3494
rect 4300 3754 4340 3794
rect 4300 3654 4340 3694
rect 4300 3554 4340 3594
rect 4300 3454 4340 3494
rect 4444 3754 4484 3794
rect 4444 3654 4484 3694
rect 4444 3554 4484 3594
rect 4444 3454 4484 3494
rect 4732 3754 4772 3794
rect 4732 3654 4772 3694
rect 4732 3554 4772 3594
rect 4732 3454 4772 3494
rect 4876 3754 4916 3794
rect 4876 3654 4916 3694
rect 4876 3554 4916 3594
rect 4876 3454 4916 3494
rect 5020 3754 5060 3794
rect 5020 3654 5060 3694
rect 5020 3554 5060 3594
rect 5020 3454 5060 3494
rect 5308 3754 5348 3794
rect 5308 3654 5348 3694
rect 5308 3554 5348 3594
rect 5308 3454 5348 3494
rect 5452 3754 5492 3794
rect 5452 3654 5492 3694
rect 5452 3554 5492 3594
rect 5452 3454 5492 3494
rect 5596 3754 5636 3794
rect 5596 3654 5636 3694
rect 5596 3554 5636 3594
rect 5596 3454 5636 3494
rect 5884 3754 5924 3794
rect 5884 3654 5924 3694
rect 5884 3554 5924 3594
rect 5884 3454 5924 3494
rect 6028 3754 6068 3794
rect 6028 3654 6068 3694
rect 6028 3554 6068 3594
rect 6028 3454 6068 3494
rect 6172 3754 6212 3794
rect 6172 3654 6212 3694
rect 6172 3554 6212 3594
rect 6172 3454 6212 3494
rect 6460 3754 6500 3794
rect 6460 3654 6500 3694
rect 6460 3554 6500 3594
rect 6460 3454 6500 3494
rect 6604 3754 6644 3794
rect 6604 3654 6644 3694
rect 6604 3554 6644 3594
rect 6604 3454 6644 3494
rect 6748 3754 6788 3794
rect 7612 3754 7652 3794
rect 6748 3654 6788 3694
rect 6748 3554 6788 3594
rect 7036 3552 7076 3704
rect 7180 3552 7220 3704
rect 7324 3552 7364 3704
rect 7612 3654 7652 3694
rect 7612 3554 7652 3594
rect 6748 3454 6788 3494
rect 7612 3454 7652 3494
rect 7756 3754 7796 3794
rect 7756 3654 7796 3694
rect 7756 3554 7796 3594
rect 7756 3454 7796 3494
rect 7900 3754 7940 3794
rect 7900 3654 7940 3694
rect 7900 3554 7940 3594
rect 7900 3454 7940 3494
rect 8188 3754 8228 3794
rect 8188 3654 8228 3694
rect 8188 3554 8228 3594
rect 8188 3454 8228 3494
rect 8332 3754 8372 3794
rect 8332 3654 8372 3694
rect 8332 3554 8372 3594
rect 8332 3454 8372 3494
rect 8476 3754 8516 3794
rect 8476 3654 8516 3694
rect 8476 3554 8516 3594
rect 8476 3454 8516 3494
rect 8764 3754 8804 3794
rect 8764 3654 8804 3694
rect 8764 3554 8804 3594
rect 8764 3454 8804 3494
rect 8908 3754 8948 3794
rect 8908 3654 8948 3694
rect 8908 3554 8948 3594
rect 8908 3454 8948 3494
rect 9052 3754 9092 3794
rect 9052 3654 9092 3694
rect 9052 3554 9092 3594
rect 9052 3454 9092 3494
rect 9340 3754 9380 3794
rect 9340 3654 9380 3694
rect 9340 3554 9380 3594
rect 9340 3454 9380 3494
rect 9484 3754 9524 3794
rect 9484 3654 9524 3694
rect 9484 3554 9524 3594
rect 9484 3454 9524 3494
rect 9628 3754 9668 3794
rect 9628 3654 9668 3694
rect 9628 3554 9668 3594
rect 9628 3454 9668 3494
rect 10204 3754 10244 3794
rect 10204 3654 10244 3694
rect 10204 3554 10244 3594
rect 10204 3454 10244 3494
rect 10348 3754 10388 3794
rect 10348 3654 10388 3694
rect 10348 3554 10388 3594
rect 10348 3454 10388 3494
rect 10492 3754 10532 3794
rect 10492 3654 10532 3694
rect 10492 3554 10532 3594
rect 10492 3454 10532 3494
rect 10780 3754 10820 3794
rect 10780 3654 10820 3694
rect 10780 3554 10820 3594
rect 10780 3454 10820 3494
rect 10924 3754 10964 3794
rect 10924 3654 10964 3694
rect 10924 3554 10964 3594
rect 10924 3454 10964 3494
rect 11068 3754 11108 3794
rect 11932 3754 11972 3794
rect 11068 3654 11108 3694
rect 11068 3554 11108 3594
rect 11356 3552 11396 3704
rect 11500 3552 11540 3704
rect 11644 3552 11684 3704
rect 11932 3654 11972 3694
rect 11932 3554 11972 3594
rect 11068 3454 11108 3494
rect 11932 3454 11972 3494
rect 12076 3754 12116 3794
rect 12076 3654 12116 3694
rect 12076 3554 12116 3594
rect 12076 3454 12116 3494
rect 12220 3754 12260 3794
rect 12220 3654 12260 3694
rect 12220 3554 12260 3594
rect 12220 3454 12260 3494
rect 12508 3754 12548 3794
rect 12508 3654 12548 3694
rect 12508 3554 12548 3594
rect 12508 3454 12548 3494
rect 12652 3754 12692 3794
rect 12652 3654 12692 3694
rect 12652 3554 12692 3594
rect 12652 3454 12692 3494
rect 12796 3754 12836 3794
rect 12796 3654 12836 3694
rect 12796 3554 12836 3594
rect 12796 3454 12836 3494
rect 13660 3754 13700 3794
rect 13660 3654 13700 3694
rect 13660 3554 13700 3594
rect 13660 3454 13700 3494
rect 13804 3754 13844 3794
rect 13804 3654 13844 3694
rect 13804 3554 13844 3594
rect 13804 3454 13844 3494
rect 13948 3754 13988 3794
rect 13948 3654 13988 3694
rect 13948 3554 13988 3594
rect 13948 3454 13988 3494
rect 14236 3754 14276 3794
rect 14236 3654 14276 3694
rect 14236 3554 14276 3594
rect 14236 3454 14276 3494
rect 14380 3754 14420 3794
rect 14380 3654 14420 3694
rect 14380 3554 14420 3594
rect 14380 3454 14420 3494
rect 14524 3754 14564 3794
rect 14524 3654 14564 3694
rect 14524 3554 14564 3594
rect 14524 3454 14564 3494
rect 14812 3754 14852 3794
rect 14812 3654 14852 3694
rect 14812 3554 14852 3594
rect 14812 3454 14852 3494
rect 14956 3754 14996 3794
rect 14956 3654 14996 3694
rect 14956 3554 14996 3594
rect 14956 3454 14996 3494
rect 15100 3754 15140 3794
rect 16540 3754 16580 3794
rect 15100 3654 15140 3694
rect 15100 3554 15140 3594
rect 15388 3552 15428 3704
rect 15532 3552 15572 3704
rect 15676 3552 15716 3704
rect 15964 3552 16004 3704
rect 16108 3552 16148 3704
rect 16252 3552 16292 3704
rect 16540 3654 16580 3694
rect 16540 3554 16580 3594
rect 15100 3454 15140 3494
rect 16540 3454 16580 3494
rect 16684 3754 16724 3794
rect 16684 3654 16724 3694
rect 16684 3554 16724 3594
rect 16684 3454 16724 3494
rect 16828 3754 16868 3794
rect 16828 3654 16868 3694
rect 16828 3554 16868 3594
rect 16828 3454 16868 3494
rect 16972 3754 17012 3794
rect 16972 3654 17012 3694
rect 16972 3554 17012 3594
rect 16972 3454 17012 3494
rect 17116 3754 17156 3794
rect 17116 3654 17156 3694
rect 17116 3554 17156 3594
rect 17116 3454 17156 3494
rect 17260 3754 17300 3794
rect 17260 3654 17300 3694
rect 17260 3554 17300 3594
rect 17260 3454 17300 3494
rect 17404 3754 17444 3794
rect 17404 3654 17444 3694
rect 17404 3554 17444 3594
rect 17404 3454 17444 3494
rect 17548 3754 17588 3794
rect 17548 3654 17588 3694
rect 17548 3554 17588 3594
rect 17548 3454 17588 3494
rect 17692 3754 17732 3794
rect 17692 3654 17732 3694
rect 17692 3554 17732 3594
rect 17692 3454 17732 3494
rect 17836 3754 17876 3794
rect 17836 3654 17876 3694
rect 17836 3554 17876 3594
rect 17836 3454 17876 3494
rect 17980 3754 18020 3794
rect 17980 3654 18020 3694
rect 17980 3554 18020 3594
rect 17980 3454 18020 3494
rect 18124 3754 18164 3794
rect 18124 3654 18164 3694
rect 18124 3554 18164 3594
rect 18124 3454 18164 3494
rect 18268 3754 18308 3794
rect 18268 3654 18308 3694
rect 18268 3554 18308 3594
rect 18268 3454 18308 3494
rect 18412 3754 18452 3794
rect 18412 3654 18452 3694
rect 18412 3554 18452 3594
rect 18412 3454 18452 3494
rect 18556 3754 18596 3794
rect 18556 3654 18596 3694
rect 18556 3554 18596 3594
rect 18556 3454 18596 3494
rect 18700 3754 18740 3794
rect 18700 3654 18740 3694
rect 18700 3554 18740 3594
rect 18700 3454 18740 3494
rect 18844 3754 18884 3794
rect 18844 3654 18884 3694
rect 18844 3554 18884 3594
rect 18844 3454 18884 3494
rect 18988 3754 19028 3794
rect 18988 3654 19028 3694
rect 18988 3554 19028 3594
rect 18988 3454 19028 3494
rect 19132 3754 19172 3794
rect 19132 3654 19172 3694
rect 19132 3554 19172 3594
rect 19132 3454 19172 3494
rect 19276 3754 19316 3794
rect 19276 3654 19316 3694
rect 19276 3554 19316 3594
rect 19276 3454 19316 3494
rect 19420 3754 19460 3794
rect 19420 3654 19460 3694
rect 19420 3554 19460 3594
rect 19420 3454 19460 3494
rect 19564 3754 19604 3794
rect 19564 3654 19604 3694
rect 19564 3554 19604 3594
rect 19564 3454 19604 3494
rect 19708 3754 19748 3794
rect 19708 3654 19748 3694
rect 19708 3554 19748 3594
rect 19708 3454 19748 3494
rect 19852 3754 19892 3794
rect 19852 3654 19892 3694
rect 19852 3554 19892 3594
rect 19852 3454 19892 3494
rect 19996 3754 20036 3794
rect 19996 3654 20036 3694
rect 19996 3554 20036 3594
rect 19996 3454 20036 3494
rect 790 3295 824 3329
rect 898 3295 932 3329
rect 1366 3295 1400 3329
rect 1474 3295 1508 3329
rect 1942 3295 1976 3329
rect 2050 3295 2084 3329
rect 2518 3295 2552 3329
rect 2626 3295 2660 3329
rect 3100 3295 3134 3329
rect 3208 3295 3242 3329
rect 4252 3295 4286 3329
rect 4360 3295 4394 3329
rect 4828 3295 4862 3329
rect 4936 3295 4970 3329
rect 5404 3295 5438 3329
rect 5512 3295 5546 3329
rect 5980 3295 6014 3329
rect 6088 3295 6122 3329
rect 6468 3294 6504 3330
rect 6752 3294 6788 3330
rect 7708 3295 7742 3329
rect 7816 3295 7850 3329
rect 8284 3295 8318 3329
rect 8392 3295 8426 3329
rect 8860 3295 8894 3329
rect 8968 3295 9002 3329
rect 9348 3294 9384 3330
rect 9632 3294 9668 3330
rect 10300 3295 10334 3329
rect 10408 3295 10442 3329
rect 10876 3295 10910 3329
rect 10984 3295 11018 3329
rect 12028 3295 12062 3329
rect 12136 3295 12170 3329
rect 12604 3295 12638 3329
rect 12712 3295 12746 3329
rect 13756 3295 13790 3329
rect 13864 3295 13898 3329
rect 14332 3295 14366 3329
rect 14440 3295 14474 3329
rect 14908 3295 14942 3329
rect 15016 3295 15050 3329
rect 16630 3295 16664 3329
rect 16738 3295 16772 3329
rect 16918 3295 16952 3329
rect 17026 3295 17060 3329
rect 17206 3295 17240 3329
rect 17314 3295 17348 3329
rect 17494 3295 17528 3329
rect 17602 3295 17636 3329
rect 17782 3295 17816 3329
rect 17890 3295 17924 3329
rect 18070 3295 18104 3329
rect 18178 3295 18212 3329
rect 18358 3295 18392 3329
rect 18466 3295 18500 3329
rect 18646 3295 18680 3329
rect 18754 3295 18788 3329
rect 18934 3295 18968 3329
rect 19042 3295 19076 3329
rect 19222 3295 19256 3329
rect 19330 3295 19364 3329
rect 19510 3295 19544 3329
rect 19618 3295 19652 3329
rect 19798 3295 19832 3329
rect 19906 3295 19940 3329
rect 790 2719 824 2753
rect 898 2719 932 2753
rect 1366 2719 1400 2753
rect 1474 2719 1508 2753
rect 1942 2719 1976 2753
rect 2050 2719 2084 2753
rect 2518 2719 2552 2753
rect 2626 2719 2660 2753
rect 3100 2719 3134 2753
rect 3208 2719 3242 2753
rect 4252 2719 4286 2753
rect 4360 2719 4394 2753
rect 4828 2719 4862 2753
rect 4936 2719 4970 2753
rect 5404 2719 5438 2753
rect 5512 2719 5546 2753
rect 5980 2719 6014 2753
rect 6088 2719 6122 2753
rect 6468 2718 6504 2754
rect 6746 2718 6782 2754
rect 7708 2719 7742 2753
rect 7816 2719 7850 2753
rect 8284 2719 8318 2753
rect 8392 2719 8426 2753
rect 8860 2719 8894 2753
rect 8968 2719 9002 2753
rect 9348 2718 9384 2754
rect 9626 2718 9662 2754
rect 10300 2719 10334 2753
rect 10408 2719 10442 2753
rect 10876 2719 10910 2753
rect 10984 2719 11018 2753
rect 12028 2719 12062 2753
rect 12136 2719 12170 2753
rect 12604 2719 12638 2753
rect 12712 2719 12746 2753
rect 13756 2719 13790 2753
rect 13864 2719 13898 2753
rect 14332 2719 14366 2753
rect 14440 2719 14474 2753
rect 14908 2719 14942 2753
rect 15016 2719 15050 2753
rect 16630 2719 16664 2753
rect 16738 2719 16772 2753
rect 16918 2719 16952 2753
rect 17026 2719 17060 2753
rect 17206 2719 17240 2753
rect 17314 2719 17348 2753
rect 17494 2719 17528 2753
rect 17602 2719 17636 2753
rect 17782 2719 17816 2753
rect 17890 2719 17924 2753
rect 18070 2719 18104 2753
rect 18178 2719 18212 2753
rect 18358 2719 18392 2753
rect 18466 2719 18500 2753
rect 18646 2719 18680 2753
rect 18754 2719 18788 2753
rect 18934 2719 18968 2753
rect 19042 2719 19076 2753
rect 19222 2719 19256 2753
rect 19330 2719 19364 2753
rect 19510 2719 19544 2753
rect 19618 2719 19652 2753
rect 19798 2719 19832 2753
rect 19906 2719 19940 2753
rect 124 2500 164 2588
rect 268 2500 308 2588
rect 412 2500 452 2588
rect 700 2574 740 2614
rect 700 2474 740 2514
rect 844 2574 884 2614
rect 844 2474 884 2514
rect 988 2574 1028 2614
rect 988 2474 1028 2514
rect 1276 2574 1316 2614
rect 1276 2474 1316 2514
rect 1420 2574 1460 2614
rect 1420 2474 1460 2514
rect 1564 2574 1604 2614
rect 1564 2474 1604 2514
rect 1852 2574 1892 2614
rect 1852 2474 1892 2514
rect 1996 2574 2036 2614
rect 1996 2474 2036 2514
rect 2140 2574 2180 2614
rect 2140 2474 2180 2514
rect 2428 2574 2468 2614
rect 2428 2474 2468 2514
rect 2572 2574 2612 2614
rect 2572 2474 2612 2514
rect 2716 2574 2756 2614
rect 2716 2474 2756 2514
rect 3004 2574 3044 2614
rect 3004 2474 3044 2514
rect 3148 2574 3188 2614
rect 3148 2474 3188 2514
rect 3292 2574 3332 2614
rect 3292 2474 3332 2514
rect 3580 2500 3620 2588
rect 3724 2500 3764 2588
rect 3868 2500 3908 2588
rect 4156 2574 4196 2614
rect 4156 2474 4196 2514
rect 4300 2574 4340 2614
rect 4300 2474 4340 2514
rect 4444 2574 4484 2614
rect 4444 2474 4484 2514
rect 4732 2574 4772 2614
rect 4732 2474 4772 2514
rect 4876 2574 4916 2614
rect 4876 2474 4916 2514
rect 5020 2574 5060 2614
rect 5020 2474 5060 2514
rect 5308 2574 5348 2614
rect 5308 2474 5348 2514
rect 5452 2574 5492 2614
rect 5452 2474 5492 2514
rect 5596 2574 5636 2614
rect 5596 2474 5636 2514
rect 5884 2574 5924 2614
rect 5884 2474 5924 2514
rect 6028 2574 6068 2614
rect 6028 2474 6068 2514
rect 6172 2574 6212 2614
rect 6172 2474 6212 2514
rect 6460 2574 6500 2614
rect 6460 2474 6500 2514
rect 6604 2574 6644 2614
rect 6604 2474 6644 2514
rect 6748 2574 6788 2614
rect 6748 2474 6788 2514
rect 7036 2500 7076 2588
rect 7180 2500 7220 2588
rect 7324 2500 7364 2588
rect 7612 2574 7652 2614
rect 7612 2474 7652 2514
rect 7756 2574 7796 2614
rect 7756 2474 7796 2514
rect 7900 2574 7940 2614
rect 7900 2474 7940 2514
rect 8188 2574 8228 2614
rect 8188 2474 8228 2514
rect 8332 2574 8372 2614
rect 8332 2474 8372 2514
rect 8476 2574 8516 2614
rect 8476 2474 8516 2514
rect 8764 2574 8804 2614
rect 8764 2474 8804 2514
rect 8908 2574 8948 2614
rect 8908 2474 8948 2514
rect 9052 2574 9092 2614
rect 9052 2474 9092 2514
rect 9340 2574 9380 2614
rect 9340 2474 9380 2514
rect 9484 2574 9524 2614
rect 9484 2474 9524 2514
rect 9628 2574 9668 2614
rect 9628 2474 9668 2514
rect 10204 2574 10244 2614
rect 10204 2474 10244 2514
rect 10348 2574 10388 2614
rect 10348 2474 10388 2514
rect 10492 2574 10532 2614
rect 10492 2474 10532 2514
rect 10780 2574 10820 2614
rect 10780 2474 10820 2514
rect 10924 2574 10964 2614
rect 10924 2474 10964 2514
rect 11068 2574 11108 2614
rect 11068 2474 11108 2514
rect 11356 2500 11396 2588
rect 11500 2500 11540 2588
rect 11644 2500 11684 2588
rect 11932 2574 11972 2614
rect 11932 2474 11972 2514
rect 12076 2574 12116 2614
rect 12076 2474 12116 2514
rect 12220 2574 12260 2614
rect 12220 2474 12260 2514
rect 12508 2574 12548 2614
rect 12508 2474 12548 2514
rect 12652 2574 12692 2614
rect 12652 2474 12692 2514
rect 12796 2574 12836 2614
rect 12796 2474 12836 2514
rect 13660 2574 13700 2614
rect 13660 2474 13700 2514
rect 13804 2574 13844 2614
rect 13804 2474 13844 2514
rect 13948 2574 13988 2614
rect 13948 2474 13988 2514
rect 14236 2574 14276 2614
rect 14236 2474 14276 2514
rect 14380 2574 14420 2614
rect 14380 2474 14420 2514
rect 14524 2574 14564 2614
rect 14524 2474 14564 2514
rect 14812 2574 14852 2614
rect 14812 2474 14852 2514
rect 14956 2574 14996 2614
rect 14956 2474 14996 2514
rect 15100 2574 15140 2614
rect 15100 2474 15140 2514
rect 15388 2500 15428 2588
rect 15532 2500 15572 2588
rect 15676 2500 15716 2588
rect 15964 2500 16004 2588
rect 16108 2500 16148 2588
rect 16252 2500 16292 2588
rect 16540 2574 16580 2614
rect 16540 2474 16580 2514
rect 16684 2574 16724 2614
rect 16684 2474 16724 2514
rect 16828 2574 16868 2614
rect 16828 2474 16868 2514
rect 16972 2574 17012 2614
rect 16972 2474 17012 2514
rect 17116 2574 17156 2614
rect 17116 2474 17156 2514
rect 17260 2574 17300 2614
rect 17260 2474 17300 2514
rect 17404 2574 17444 2614
rect 17404 2474 17444 2514
rect 17548 2574 17588 2614
rect 17548 2474 17588 2514
rect 17692 2574 17732 2614
rect 17692 2474 17732 2514
rect 17836 2574 17876 2614
rect 17836 2474 17876 2514
rect 17980 2574 18020 2614
rect 17980 2474 18020 2514
rect 18124 2574 18164 2614
rect 18124 2474 18164 2514
rect 18268 2574 18308 2614
rect 18268 2474 18308 2514
rect 18412 2574 18452 2614
rect 18412 2474 18452 2514
rect 18556 2574 18596 2614
rect 18556 2474 18596 2514
rect 18700 2574 18740 2614
rect 18700 2474 18740 2514
rect 18844 2574 18884 2614
rect 18844 2474 18884 2514
rect 18988 2574 19028 2614
rect 18988 2474 19028 2514
rect 19132 2574 19172 2614
rect 19132 2474 19172 2514
rect 19276 2574 19316 2614
rect 19276 2474 19316 2514
rect 19420 2574 19460 2614
rect 19420 2474 19460 2514
rect 19564 2574 19604 2614
rect 19564 2474 19604 2514
rect 19708 2574 19748 2614
rect 19708 2474 19748 2514
rect 19852 2574 19892 2614
rect 19852 2474 19892 2514
rect 19996 2574 20036 2614
rect 19996 2474 20036 2514
rect 124 1444 164 1532
rect 268 1444 308 1532
rect 412 1444 452 1532
rect 700 1518 740 1558
rect 700 1418 740 1458
rect 844 1518 884 1558
rect 844 1418 884 1458
rect 988 1518 1028 1558
rect 988 1418 1028 1458
rect 1276 1518 1316 1558
rect 1276 1418 1316 1458
rect 1420 1518 1460 1558
rect 1420 1418 1460 1458
rect 1564 1518 1604 1558
rect 1564 1418 1604 1458
rect 1852 1518 1892 1558
rect 1852 1418 1892 1458
rect 1996 1518 2036 1558
rect 1996 1418 2036 1458
rect 2140 1518 2180 1558
rect 2140 1418 2180 1458
rect 3004 1518 3044 1558
rect 3004 1418 3044 1458
rect 3148 1518 3188 1558
rect 3148 1418 3188 1458
rect 3292 1518 3332 1558
rect 3292 1418 3332 1458
rect 3580 1518 3620 1558
rect 3580 1418 3620 1458
rect 3724 1518 3764 1558
rect 3724 1418 3764 1458
rect 3868 1518 3908 1558
rect 3868 1418 3908 1458
rect 4156 1518 4196 1558
rect 4156 1418 4196 1458
rect 4300 1518 4340 1558
rect 4300 1418 4340 1458
rect 4444 1518 4484 1558
rect 4444 1418 4484 1458
rect 4732 1444 4772 1532
rect 4876 1444 4916 1532
rect 5020 1444 5060 1532
rect 5308 1444 5348 1532
rect 5452 1444 5492 1532
rect 5596 1444 5636 1532
rect 5884 1518 5924 1558
rect 5884 1418 5924 1458
rect 6028 1518 6068 1558
rect 6028 1418 6068 1458
rect 6172 1518 6212 1558
rect 6172 1418 6212 1458
rect 6460 1518 6500 1558
rect 6460 1418 6500 1458
rect 6604 1518 6644 1558
rect 6604 1418 6644 1458
rect 6748 1518 6788 1558
rect 6748 1418 6788 1458
rect 7036 1518 7076 1558
rect 7036 1418 7076 1458
rect 7180 1518 7220 1558
rect 7180 1418 7220 1458
rect 7324 1518 7364 1558
rect 7324 1418 7364 1458
rect 7612 1518 7652 1558
rect 7612 1418 7652 1458
rect 7756 1518 7796 1558
rect 7756 1418 7796 1458
rect 7900 1518 7940 1558
rect 7900 1418 7940 1458
rect 8188 1518 8228 1558
rect 8188 1418 8228 1458
rect 8332 1518 8372 1558
rect 8332 1418 8372 1458
rect 8476 1518 8516 1558
rect 8476 1418 8516 1458
rect 8764 1444 8804 1532
rect 8908 1444 8948 1532
rect 9052 1444 9092 1532
rect 9340 1518 9380 1558
rect 9340 1418 9380 1458
rect 9484 1518 9524 1558
rect 9484 1418 9524 1458
rect 9628 1518 9668 1558
rect 9628 1418 9668 1458
rect 9916 1518 9956 1558
rect 9916 1418 9956 1458
rect 10060 1518 10100 1558
rect 10060 1418 10100 1458
rect 10204 1518 10244 1558
rect 10204 1418 10244 1458
rect 10492 1518 10532 1558
rect 10492 1418 10532 1458
rect 10636 1518 10676 1558
rect 10636 1418 10676 1458
rect 10780 1518 10820 1558
rect 10780 1418 10820 1458
rect 11068 1518 11108 1558
rect 11068 1418 11108 1458
rect 11212 1518 11252 1558
rect 11212 1418 11252 1458
rect 11356 1518 11396 1558
rect 11356 1418 11396 1458
rect 11932 1518 11972 1558
rect 11932 1418 11972 1458
rect 12076 1518 12116 1558
rect 12076 1418 12116 1458
rect 12220 1518 12260 1558
rect 12220 1418 12260 1458
rect 12508 1518 12548 1558
rect 12508 1418 12548 1458
rect 12652 1518 12692 1558
rect 12652 1418 12692 1458
rect 12796 1518 12836 1558
rect 12796 1418 12836 1458
rect 13084 1518 13124 1558
rect 13084 1418 13124 1458
rect 13228 1518 13268 1558
rect 13228 1418 13268 1458
rect 13372 1518 13412 1558
rect 13372 1418 13412 1458
rect 13660 1518 13700 1558
rect 13660 1418 13700 1458
rect 13804 1518 13844 1558
rect 13804 1418 13844 1458
rect 13948 1518 13988 1558
rect 13948 1418 13988 1458
rect 14236 1444 14276 1532
rect 14380 1444 14420 1532
rect 14524 1444 14564 1532
rect 14812 1518 14852 1558
rect 14812 1418 14852 1458
rect 14956 1518 14996 1558
rect 14956 1418 14996 1458
rect 15100 1518 15140 1558
rect 15100 1418 15140 1458
rect 15388 1518 15428 1558
rect 15388 1418 15428 1458
rect 15532 1518 15572 1558
rect 15532 1418 15572 1458
rect 15676 1518 15716 1558
rect 15676 1418 15716 1458
rect 15964 1518 16004 1558
rect 15964 1418 16004 1458
rect 16108 1518 16148 1558
rect 16108 1418 16148 1458
rect 16252 1518 16292 1558
rect 16252 1418 16292 1458
rect 16396 1518 16436 1558
rect 16396 1418 16436 1458
rect 16540 1518 16580 1558
rect 16540 1418 16580 1458
rect 16828 1444 16868 1532
rect 16972 1444 17012 1532
rect 17116 1444 17156 1532
rect 17404 1518 17444 1558
rect 17404 1418 17444 1458
rect 17548 1518 17588 1558
rect 17548 1418 17588 1458
rect 17692 1518 17732 1558
rect 17692 1418 17732 1458
rect 17836 1518 17876 1558
rect 17836 1418 17876 1458
rect 17980 1518 18020 1558
rect 17980 1418 18020 1458
rect 18124 1518 18164 1558
rect 18124 1418 18164 1458
rect 18268 1518 18308 1558
rect 18268 1418 18308 1458
rect 18412 1518 18452 1558
rect 18412 1418 18452 1458
rect 18556 1518 18596 1558
rect 18556 1418 18596 1458
rect 18700 1518 18740 1558
rect 18700 1418 18740 1458
rect 18844 1518 18884 1558
rect 18844 1418 18884 1458
rect 18988 1518 19028 1558
rect 18988 1418 19028 1458
rect 19132 1518 19172 1558
rect 19132 1418 19172 1458
rect 19276 1518 19316 1558
rect 19276 1418 19316 1458
rect 19420 1518 19460 1558
rect 19420 1418 19460 1458
rect 19564 1518 19604 1558
rect 19564 1418 19604 1458
rect 19708 1518 19748 1558
rect 19708 1418 19748 1458
rect 19852 1518 19892 1558
rect 19852 1418 19892 1458
rect 19996 1518 20036 1558
rect 19996 1418 20036 1458
rect 20140 1518 20180 1558
rect 20140 1418 20180 1458
rect 20284 1518 20324 1558
rect 20284 1418 20324 1458
rect 20428 1518 20468 1558
rect 20428 1418 20468 1458
rect 20572 1518 20612 1558
rect 20572 1418 20612 1458
rect 20716 1518 20756 1558
rect 20716 1418 20756 1458
rect 20860 1518 20900 1558
rect 20860 1418 20900 1458
rect 796 1279 830 1313
rect 904 1279 938 1313
rect 1372 1279 1406 1313
rect 1480 1279 1514 1313
rect 1948 1279 1982 1313
rect 2056 1279 2090 1313
rect 3100 1279 3134 1313
rect 3208 1279 3242 1313
rect 3676 1279 3710 1313
rect 3784 1279 3818 1313
rect 4252 1279 4286 1313
rect 4360 1279 4394 1313
rect 5980 1279 6014 1313
rect 6088 1279 6122 1313
rect 6556 1279 6590 1313
rect 6664 1279 6698 1313
rect 7132 1279 7166 1313
rect 7240 1279 7274 1313
rect 7708 1279 7742 1313
rect 7816 1279 7850 1313
rect 8196 1278 8232 1314
rect 8474 1278 8510 1314
rect 9436 1279 9470 1313
rect 9544 1279 9578 1313
rect 10012 1279 10046 1313
rect 10120 1279 10154 1313
rect 10588 1279 10622 1313
rect 10696 1279 10730 1313
rect 11076 1278 11112 1314
rect 11354 1278 11390 1314
rect 12028 1279 12062 1313
rect 12136 1279 12170 1313
rect 12604 1279 12638 1313
rect 12712 1279 12746 1313
rect 13180 1279 13214 1313
rect 13288 1279 13322 1313
rect 13756 1279 13790 1313
rect 13864 1279 13898 1313
rect 14908 1279 14942 1313
rect 15016 1279 15050 1313
rect 15478 1279 15512 1313
rect 15586 1279 15620 1313
rect 16060 1279 16094 1313
rect 16168 1279 16202 1313
rect 16348 1279 16382 1313
rect 16456 1279 16490 1313
rect 17500 1279 17534 1313
rect 17608 1279 17642 1313
rect 17788 1279 17822 1313
rect 17896 1279 17930 1313
rect 18076 1279 18110 1313
rect 18184 1279 18218 1313
rect 18364 1279 18398 1313
rect 18472 1279 18506 1313
rect 18652 1279 18686 1313
rect 18760 1279 18794 1313
rect 18940 1279 18974 1313
rect 19048 1279 19082 1313
rect 19228 1279 19262 1313
rect 19336 1279 19370 1313
rect 19516 1279 19550 1313
rect 19624 1279 19658 1313
rect 19804 1279 19838 1313
rect 19912 1279 19946 1313
rect 20092 1279 20126 1313
rect 20200 1279 20234 1313
rect 20380 1279 20414 1313
rect 20488 1279 20522 1313
rect 20668 1279 20702 1313
rect 20776 1279 20810 1313
rect 796 703 830 737
rect 904 703 938 737
rect 1372 703 1406 737
rect 1480 703 1514 737
rect 1948 703 1982 737
rect 2056 703 2090 737
rect 3100 703 3134 737
rect 3208 703 3242 737
rect 3676 703 3710 737
rect 3784 703 3818 737
rect 4252 703 4286 737
rect 4360 703 4394 737
rect 5980 703 6014 737
rect 6088 703 6122 737
rect 6556 703 6590 737
rect 6664 703 6698 737
rect 7132 703 7166 737
rect 7240 703 7274 737
rect 7708 703 7742 737
rect 7816 703 7850 737
rect 8196 702 8232 738
rect 8480 702 8516 738
rect 9436 703 9470 737
rect 9544 703 9578 737
rect 10012 703 10046 737
rect 10120 703 10154 737
rect 10588 703 10622 737
rect 10696 703 10730 737
rect 11076 702 11112 738
rect 11360 702 11396 738
rect 12028 703 12062 737
rect 12136 703 12170 737
rect 12604 703 12638 737
rect 12712 703 12746 737
rect 13180 703 13214 737
rect 13288 703 13322 737
rect 13756 703 13790 737
rect 13864 703 13898 737
rect 14908 703 14942 737
rect 15016 703 15050 737
rect 15478 703 15512 737
rect 15586 703 15620 737
rect 16060 703 16094 737
rect 16168 703 16202 737
rect 16348 703 16382 737
rect 16456 703 16490 737
rect 17500 703 17534 737
rect 17608 703 17642 737
rect 17788 703 17822 737
rect 17896 703 17930 737
rect 18076 703 18110 737
rect 18184 703 18218 737
rect 18364 703 18398 737
rect 18472 703 18506 737
rect 18652 703 18686 737
rect 18760 703 18794 737
rect 18940 703 18974 737
rect 19048 703 19082 737
rect 19228 703 19262 737
rect 19336 703 19370 737
rect 19516 703 19550 737
rect 19624 703 19658 737
rect 19804 703 19838 737
rect 19912 703 19946 737
rect 20092 703 20126 737
rect 20200 703 20234 737
rect 20380 703 20414 737
rect 20488 703 20522 737
rect 20668 703 20702 737
rect 20776 703 20810 737
rect 700 538 740 578
rect 124 328 164 480
rect 268 328 308 480
rect 412 328 452 480
rect 700 438 740 478
rect 700 338 740 378
rect 700 238 740 278
rect 844 538 884 578
rect 844 438 884 478
rect 844 338 884 378
rect 844 238 884 278
rect 988 538 1028 578
rect 988 438 1028 478
rect 988 338 1028 378
rect 988 238 1028 278
rect 1276 538 1316 578
rect 1276 438 1316 478
rect 1276 338 1316 378
rect 1276 238 1316 278
rect 1420 538 1460 578
rect 1420 438 1460 478
rect 1420 338 1460 378
rect 1420 238 1460 278
rect 1564 538 1604 578
rect 1564 438 1604 478
rect 1564 338 1604 378
rect 1564 238 1604 278
rect 1852 538 1892 578
rect 1852 438 1892 478
rect 1852 338 1892 378
rect 1852 238 1892 278
rect 1996 538 2036 578
rect 1996 438 2036 478
rect 1996 338 2036 378
rect 1996 238 2036 278
rect 2140 538 2180 578
rect 2140 438 2180 478
rect 2140 338 2180 378
rect 2140 238 2180 278
rect 3004 538 3044 578
rect 3004 438 3044 478
rect 3004 338 3044 378
rect 3004 238 3044 278
rect 3148 538 3188 578
rect 3148 438 3188 478
rect 3148 338 3188 378
rect 3148 238 3188 278
rect 3292 538 3332 578
rect 3292 438 3332 478
rect 3292 338 3332 378
rect 3292 238 3332 278
rect 3580 538 3620 578
rect 3580 438 3620 478
rect 3580 338 3620 378
rect 3580 238 3620 278
rect 3724 538 3764 578
rect 3724 438 3764 478
rect 3724 338 3764 378
rect 3724 238 3764 278
rect 3868 538 3908 578
rect 3868 438 3908 478
rect 3868 338 3908 378
rect 3868 238 3908 278
rect 4156 538 4196 578
rect 4156 438 4196 478
rect 4156 338 4196 378
rect 4156 238 4196 278
rect 4300 538 4340 578
rect 4300 438 4340 478
rect 4300 338 4340 378
rect 4300 238 4340 278
rect 4444 538 4484 578
rect 5884 538 5924 578
rect 4444 438 4484 478
rect 4444 338 4484 378
rect 4732 328 4772 480
rect 4876 328 4916 480
rect 5020 328 5060 480
rect 5308 328 5348 480
rect 5452 328 5492 480
rect 5596 328 5636 480
rect 5884 438 5924 478
rect 5884 338 5924 378
rect 4444 238 4484 278
rect 5884 238 5924 278
rect 6028 538 6068 578
rect 6028 438 6068 478
rect 6028 338 6068 378
rect 6028 238 6068 278
rect 6172 538 6212 578
rect 6172 438 6212 478
rect 6172 338 6212 378
rect 6172 238 6212 278
rect 6460 538 6500 578
rect 6460 438 6500 478
rect 6460 338 6500 378
rect 6460 238 6500 278
rect 6604 538 6644 578
rect 6604 438 6644 478
rect 6604 338 6644 378
rect 6604 238 6644 278
rect 6748 538 6788 578
rect 6748 438 6788 478
rect 6748 338 6788 378
rect 6748 238 6788 278
rect 7036 538 7076 578
rect 7036 438 7076 478
rect 7036 338 7076 378
rect 7036 238 7076 278
rect 7180 538 7220 578
rect 7180 438 7220 478
rect 7180 338 7220 378
rect 7180 238 7220 278
rect 7324 538 7364 578
rect 7324 438 7364 478
rect 7324 338 7364 378
rect 7324 238 7364 278
rect 7612 538 7652 578
rect 7612 438 7652 478
rect 7612 338 7652 378
rect 7612 238 7652 278
rect 7756 538 7796 578
rect 7756 438 7796 478
rect 7756 338 7796 378
rect 7756 238 7796 278
rect 7900 538 7940 578
rect 7900 438 7940 478
rect 7900 338 7940 378
rect 7900 238 7940 278
rect 8188 538 8228 578
rect 8188 438 8228 478
rect 8188 338 8228 378
rect 8188 238 8228 278
rect 8332 538 8372 578
rect 8332 438 8372 478
rect 8332 338 8372 378
rect 8332 238 8372 278
rect 8476 538 8516 578
rect 9340 538 9380 578
rect 8476 438 8516 478
rect 8476 338 8516 378
rect 8764 328 8804 480
rect 8908 328 8948 480
rect 9052 328 9092 480
rect 9340 438 9380 478
rect 9340 338 9380 378
rect 8476 238 8516 278
rect 9340 238 9380 278
rect 9484 538 9524 578
rect 9484 438 9524 478
rect 9484 338 9524 378
rect 9484 238 9524 278
rect 9628 538 9668 578
rect 9628 438 9668 478
rect 9628 338 9668 378
rect 9628 238 9668 278
rect 9916 538 9956 578
rect 9916 438 9956 478
rect 9916 338 9956 378
rect 9916 238 9956 278
rect 10060 538 10100 578
rect 10060 438 10100 478
rect 10060 338 10100 378
rect 10060 238 10100 278
rect 10204 538 10244 578
rect 10204 438 10244 478
rect 10204 338 10244 378
rect 10204 238 10244 278
rect 10492 538 10532 578
rect 10492 438 10532 478
rect 10492 338 10532 378
rect 10492 238 10532 278
rect 10636 538 10676 578
rect 10636 438 10676 478
rect 10636 338 10676 378
rect 10636 238 10676 278
rect 10780 538 10820 578
rect 10780 438 10820 478
rect 10780 338 10820 378
rect 10780 238 10820 278
rect 11068 538 11108 578
rect 11068 438 11108 478
rect 11068 338 11108 378
rect 11068 238 11108 278
rect 11212 538 11252 578
rect 11212 438 11252 478
rect 11212 338 11252 378
rect 11212 238 11252 278
rect 11356 538 11396 578
rect 11356 438 11396 478
rect 11356 338 11396 378
rect 11356 238 11396 278
rect 11932 538 11972 578
rect 11932 438 11972 478
rect 11932 338 11972 378
rect 11932 238 11972 278
rect 12076 538 12116 578
rect 12076 438 12116 478
rect 12076 338 12116 378
rect 12076 238 12116 278
rect 12220 538 12260 578
rect 12220 438 12260 478
rect 12220 338 12260 378
rect 12220 238 12260 278
rect 12508 538 12548 578
rect 12508 438 12548 478
rect 12508 338 12548 378
rect 12508 238 12548 278
rect 12652 538 12692 578
rect 12652 438 12692 478
rect 12652 338 12692 378
rect 12652 238 12692 278
rect 12796 538 12836 578
rect 12796 438 12836 478
rect 12796 338 12836 378
rect 12796 238 12836 278
rect 13084 538 13124 578
rect 13084 438 13124 478
rect 13084 338 13124 378
rect 13084 238 13124 278
rect 13228 538 13268 578
rect 13228 438 13268 478
rect 13228 338 13268 378
rect 13228 238 13268 278
rect 13372 538 13412 578
rect 13372 438 13412 478
rect 13372 338 13412 378
rect 13372 238 13412 278
rect 13660 538 13700 578
rect 13660 438 13700 478
rect 13660 338 13700 378
rect 13660 238 13700 278
rect 13804 538 13844 578
rect 13804 438 13844 478
rect 13804 338 13844 378
rect 13804 238 13844 278
rect 13948 538 13988 578
rect 14812 538 14852 578
rect 13948 438 13988 478
rect 13948 338 13988 378
rect 14236 328 14276 480
rect 14380 328 14420 480
rect 14524 328 14564 480
rect 14812 438 14852 478
rect 14812 338 14852 378
rect 13948 238 13988 278
rect 14812 238 14852 278
rect 14956 538 14996 578
rect 14956 438 14996 478
rect 14956 338 14996 378
rect 14956 238 14996 278
rect 15100 538 15140 578
rect 15100 438 15140 478
rect 15100 338 15140 378
rect 15100 238 15140 278
rect 15388 538 15428 578
rect 15388 438 15428 478
rect 15388 338 15428 378
rect 15388 238 15428 278
rect 15532 538 15572 578
rect 15532 438 15572 478
rect 15532 338 15572 378
rect 15532 238 15572 278
rect 15676 538 15716 578
rect 15676 438 15716 478
rect 15676 338 15716 378
rect 15676 238 15716 278
rect 15964 538 16004 578
rect 15964 438 16004 478
rect 15964 338 16004 378
rect 15964 238 16004 278
rect 16108 538 16148 578
rect 16108 438 16148 478
rect 16108 338 16148 378
rect 16108 238 16148 278
rect 16252 538 16292 578
rect 16252 438 16292 478
rect 16252 338 16292 378
rect 16252 238 16292 278
rect 16396 538 16436 578
rect 16396 438 16436 478
rect 16396 338 16436 378
rect 16396 238 16436 278
rect 16540 538 16580 578
rect 17404 538 17444 578
rect 16540 438 16580 478
rect 16540 338 16580 378
rect 16828 328 16868 480
rect 16972 328 17012 480
rect 17116 328 17156 480
rect 17404 438 17444 478
rect 17404 338 17444 378
rect 16540 238 16580 278
rect 17404 238 17444 278
rect 17548 538 17588 578
rect 17548 438 17588 478
rect 17548 338 17588 378
rect 17548 238 17588 278
rect 17692 538 17732 578
rect 17692 438 17732 478
rect 17692 338 17732 378
rect 17692 238 17732 278
rect 17836 538 17876 578
rect 17836 438 17876 478
rect 17836 338 17876 378
rect 17836 238 17876 278
rect 17980 538 18020 578
rect 17980 438 18020 478
rect 17980 338 18020 378
rect 17980 238 18020 278
rect 18124 538 18164 578
rect 18124 438 18164 478
rect 18124 338 18164 378
rect 18124 238 18164 278
rect 18268 538 18308 578
rect 18268 438 18308 478
rect 18268 338 18308 378
rect 18268 238 18308 278
rect 18412 538 18452 578
rect 18412 438 18452 478
rect 18412 338 18452 378
rect 18412 238 18452 278
rect 18556 538 18596 578
rect 18556 438 18596 478
rect 18556 338 18596 378
rect 18556 238 18596 278
rect 18700 538 18740 578
rect 18700 438 18740 478
rect 18700 338 18740 378
rect 18700 238 18740 278
rect 18844 538 18884 578
rect 18844 438 18884 478
rect 18844 338 18884 378
rect 18844 238 18884 278
rect 18988 538 19028 578
rect 18988 438 19028 478
rect 18988 338 19028 378
rect 18988 238 19028 278
rect 19132 538 19172 578
rect 19132 438 19172 478
rect 19132 338 19172 378
rect 19132 238 19172 278
rect 19276 538 19316 578
rect 19276 438 19316 478
rect 19276 338 19316 378
rect 19276 238 19316 278
rect 19420 538 19460 578
rect 19420 438 19460 478
rect 19420 338 19460 378
rect 19420 238 19460 278
rect 19564 538 19604 578
rect 19564 438 19604 478
rect 19564 338 19604 378
rect 19564 238 19604 278
rect 19708 538 19748 578
rect 19708 438 19748 478
rect 19708 338 19748 378
rect 19708 238 19748 278
rect 19852 538 19892 578
rect 19852 438 19892 478
rect 19852 338 19892 378
rect 19852 238 19892 278
rect 19996 538 20036 578
rect 19996 438 20036 478
rect 19996 338 20036 378
rect 19996 238 20036 278
rect 20140 538 20180 578
rect 20140 438 20180 478
rect 20140 338 20180 378
rect 20140 238 20180 278
rect 20284 538 20324 578
rect 20284 438 20324 478
rect 20284 338 20324 378
rect 20284 238 20324 278
rect 20428 538 20468 578
rect 20428 438 20468 478
rect 20428 338 20468 378
rect 20428 238 20468 278
rect 20572 538 20612 578
rect 20572 438 20612 478
rect 20572 338 20612 378
rect 20572 238 20612 278
rect 20716 538 20756 578
rect 20716 438 20756 478
rect 20716 338 20756 378
rect 20716 238 20756 278
rect 20860 538 20900 578
rect 20860 438 20900 478
rect 20860 338 20900 378
rect 20860 238 20900 278
<< metal1 >>
rect 114 4064 174 4072
rect 402 4064 462 4072
rect 690 4064 750 4072
rect 978 4064 1038 4072
rect 1266 4064 1326 4072
rect 1554 4064 1614 4072
rect 1842 4064 1902 4072
rect 2130 4064 2190 4072
rect 2418 4064 2478 4072
rect 2706 4064 2766 4072
rect 2994 4064 3054 4072
rect 3282 4064 3342 4072
rect 3570 4064 3630 4072
rect 3858 4064 3918 4072
rect 4146 4064 4206 4072
rect 4434 4064 4494 4072
rect 4722 4064 4782 4072
rect 5010 4064 5070 4072
rect 5298 4064 5358 4072
rect 5586 4064 5646 4072
rect 7026 4064 7086 4072
rect 7314 4064 7374 4072
rect 7602 4064 7662 4072
rect 7890 4064 7950 4072
rect 8178 4064 8238 4072
rect 8466 4064 8526 4072
rect 10194 4064 10254 4072
rect 10482 4064 10542 4072
rect 10770 4064 10830 4072
rect 11058 4064 11118 4072
rect 11346 4064 11406 4072
rect 11634 4064 11694 4072
rect 11922 4064 11982 4072
rect 12210 4064 12270 4072
rect 14226 4064 14286 4072
rect 14514 4064 14574 4072
rect 14802 4064 14862 4072
rect 15090 4064 15150 4072
rect 15378 4064 15438 4072
rect 15666 4064 15726 4072
rect 15954 4064 16014 4072
rect 16242 4064 16302 4072
rect 16530 4064 16590 4072
rect 16818 4064 16878 4072
rect 17106 4064 17166 4072
rect 17394 4064 17454 4072
rect 17682 4064 17742 4072
rect 17970 4064 18030 4072
rect 18258 4064 18318 4072
rect 18546 4064 18606 4072
rect 18834 4064 18894 4072
rect 19122 4064 19182 4072
rect 19410 4064 19470 4072
rect 19698 4064 19758 4072
rect 19986 4064 20046 4072
rect 112 4058 176 4064
rect 112 4006 118 4058
rect 170 4006 176 4058
rect 112 4000 176 4006
rect 400 4058 464 4064
rect 400 4006 406 4058
rect 458 4006 464 4058
rect 400 4000 464 4006
rect 688 4058 752 4064
rect 688 4006 694 4058
rect 746 4006 752 4058
rect 688 4000 752 4006
rect 976 4058 1040 4064
rect 976 4006 982 4058
rect 1034 4006 1040 4058
rect 976 4000 1040 4006
rect 1264 4058 1328 4064
rect 1264 4006 1270 4058
rect 1322 4006 1328 4058
rect 1264 4000 1328 4006
rect 1552 4058 1616 4064
rect 1552 4006 1558 4058
rect 1610 4006 1616 4058
rect 1552 4000 1616 4006
rect 1840 4058 1904 4064
rect 1840 4006 1846 4058
rect 1898 4006 1904 4058
rect 1840 4000 1904 4006
rect 2128 4058 2192 4064
rect 2128 4006 2134 4058
rect 2186 4006 2192 4058
rect 2128 4000 2192 4006
rect 2416 4058 2480 4064
rect 2416 4006 2422 4058
rect 2474 4006 2480 4058
rect 2416 4000 2480 4006
rect 2704 4058 2768 4064
rect 2704 4006 2710 4058
rect 2762 4006 2768 4058
rect 2704 4000 2768 4006
rect 2992 4058 3056 4064
rect 2992 4006 2998 4058
rect 3050 4006 3056 4058
rect 2992 4000 3056 4006
rect 3280 4058 3344 4064
rect 3280 4006 3286 4058
rect 3338 4006 3344 4058
rect 3280 4000 3344 4006
rect 3568 4058 3632 4064
rect 3568 4006 3574 4058
rect 3626 4006 3632 4058
rect 3568 4000 3632 4006
rect 3856 4058 3920 4064
rect 3856 4006 3862 4058
rect 3914 4006 3920 4058
rect 3856 4000 3920 4006
rect 4144 4058 4208 4064
rect 4144 4006 4150 4058
rect 4202 4006 4208 4058
rect 4144 4000 4208 4006
rect 4432 4058 4496 4064
rect 4432 4006 4438 4058
rect 4490 4006 4496 4058
rect 4432 4000 4496 4006
rect 4720 4058 4784 4064
rect 4720 4006 4726 4058
rect 4778 4006 4784 4058
rect 4720 4000 4784 4006
rect 5008 4058 5072 4064
rect 5008 4006 5014 4058
rect 5066 4006 5072 4058
rect 5008 4000 5072 4006
rect 5296 4058 5360 4064
rect 5296 4006 5302 4058
rect 5354 4006 5360 4058
rect 5296 4000 5360 4006
rect 5584 4058 5648 4064
rect 5584 4006 5590 4058
rect 5642 4006 5648 4058
rect 5584 4000 5648 4006
rect 6448 4058 6512 4064
rect 6448 4006 6454 4058
rect 6506 4006 6512 4058
rect 6448 4000 6512 4006
rect 7024 4058 7088 4064
rect 7024 4006 7030 4058
rect 7082 4006 7088 4058
rect 7024 4000 7088 4006
rect 7312 4058 7376 4064
rect 7312 4006 7318 4058
rect 7370 4006 7376 4058
rect 7312 4000 7376 4006
rect 7600 4058 7664 4064
rect 7600 4006 7606 4058
rect 7658 4006 7664 4058
rect 7600 4000 7664 4006
rect 7888 4058 7952 4064
rect 7888 4006 7894 4058
rect 7946 4006 7952 4058
rect 7888 4000 7952 4006
rect 8176 4058 8240 4064
rect 8176 4006 8182 4058
rect 8234 4006 8240 4058
rect 8176 4000 8240 4006
rect 8464 4058 8528 4064
rect 8464 4006 8470 4058
rect 8522 4006 8528 4058
rect 8464 4000 8528 4006
rect 9328 4058 9392 4064
rect 9328 4006 9334 4058
rect 9386 4006 9392 4058
rect 9328 4000 9392 4006
rect 10192 4058 10256 4064
rect 10192 4006 10198 4058
rect 10250 4006 10256 4058
rect 10192 4000 10256 4006
rect 10480 4058 10544 4064
rect 10480 4006 10486 4058
rect 10538 4006 10544 4058
rect 10480 4000 10544 4006
rect 10768 4058 10832 4064
rect 10768 4006 10774 4058
rect 10826 4006 10832 4058
rect 10768 4000 10832 4006
rect 11056 4058 11120 4064
rect 11056 4006 11062 4058
rect 11114 4006 11120 4058
rect 11056 4000 11120 4006
rect 11344 4058 11408 4064
rect 11344 4006 11350 4058
rect 11402 4006 11408 4058
rect 11344 4000 11408 4006
rect 11632 4058 11696 4064
rect 11632 4006 11638 4058
rect 11690 4006 11696 4058
rect 11632 4000 11696 4006
rect 11920 4058 11984 4064
rect 11920 4006 11926 4058
rect 11978 4006 11984 4058
rect 11920 4000 11984 4006
rect 12208 4058 12272 4064
rect 12208 4006 12214 4058
rect 12266 4006 12272 4058
rect 12208 4000 12272 4006
rect 14224 4058 14288 4064
rect 14224 4006 14230 4058
rect 14282 4006 14288 4058
rect 14224 4000 14288 4006
rect 14512 4058 14576 4064
rect 14512 4006 14518 4058
rect 14570 4006 14576 4058
rect 14512 4000 14576 4006
rect 14800 4058 14864 4064
rect 14800 4006 14806 4058
rect 14858 4006 14864 4058
rect 14800 4000 14864 4006
rect 15088 4058 15152 4064
rect 15088 4006 15094 4058
rect 15146 4006 15152 4058
rect 15088 4000 15152 4006
rect 15376 4058 15440 4064
rect 15376 4006 15382 4058
rect 15434 4006 15440 4058
rect 15376 4000 15440 4006
rect 15664 4058 15728 4064
rect 15664 4006 15670 4058
rect 15722 4006 15728 4058
rect 15664 4000 15728 4006
rect 15952 4058 16016 4064
rect 15952 4006 15958 4058
rect 16010 4006 16016 4058
rect 15952 4000 16016 4006
rect 16240 4058 16304 4064
rect 16240 4006 16246 4058
rect 16298 4006 16304 4058
rect 16240 4000 16304 4006
rect 16528 4058 16592 4064
rect 16528 4006 16534 4058
rect 16586 4006 16592 4058
rect 16528 4000 16592 4006
rect 16816 4058 16880 4064
rect 16816 4006 16822 4058
rect 16874 4006 16880 4058
rect 16816 4000 16880 4006
rect 17104 4058 17168 4064
rect 17104 4006 17110 4058
rect 17162 4006 17168 4058
rect 17104 4000 17168 4006
rect 17392 4058 17456 4064
rect 17392 4006 17398 4058
rect 17450 4006 17456 4058
rect 17392 4000 17456 4006
rect 17680 4058 17744 4064
rect 17680 4006 17686 4058
rect 17738 4006 17744 4058
rect 17680 4000 17744 4006
rect 17968 4058 18032 4064
rect 17968 4006 17974 4058
rect 18026 4006 18032 4058
rect 17968 4000 18032 4006
rect 18256 4058 18320 4064
rect 18256 4006 18262 4058
rect 18314 4006 18320 4058
rect 18256 4000 18320 4006
rect 18544 4058 18608 4064
rect 18544 4006 18550 4058
rect 18602 4006 18608 4058
rect 18544 4000 18608 4006
rect 18832 4058 18896 4064
rect 18832 4006 18838 4058
rect 18890 4006 18896 4058
rect 18832 4000 18896 4006
rect 19120 4058 19184 4064
rect 19120 4006 19126 4058
rect 19178 4006 19184 4058
rect 19120 4000 19184 4006
rect 19408 4058 19472 4064
rect 19408 4006 19414 4058
rect 19466 4006 19472 4058
rect 19408 4000 19472 4006
rect 19696 4058 19760 4064
rect 19696 4006 19702 4058
rect 19754 4006 19760 4058
rect 19696 4000 19760 4006
rect 19984 4058 20048 4064
rect 19984 4006 19990 4058
rect 20042 4006 20048 4058
rect 19984 4000 20048 4006
rect 114 3704 174 4000
rect 114 3552 124 3704
rect 164 3552 174 3704
rect 258 3704 318 3844
rect 258 3632 268 3704
rect 256 3626 268 3632
rect 308 3632 318 3704
rect 402 3704 462 4000
rect 308 3626 320 3632
rect 256 3574 262 3626
rect 314 3574 320 3626
rect 256 3568 268 3574
rect 114 3528 174 3552
rect 258 3552 268 3568
rect 308 3568 320 3574
rect 308 3552 318 3568
rect 258 3528 318 3552
rect 402 3552 412 3704
rect 452 3552 462 3704
rect 402 3528 462 3552
rect 690 3794 750 4000
rect 690 3754 700 3794
rect 740 3754 750 3794
rect 690 3694 750 3754
rect 690 3654 700 3694
rect 740 3654 750 3694
rect 690 3594 750 3654
rect 834 3794 894 3844
rect 834 3754 844 3794
rect 884 3754 894 3794
rect 834 3694 894 3754
rect 834 3654 844 3694
rect 884 3654 894 3694
rect 834 3632 894 3654
rect 978 3794 1038 4000
rect 978 3754 988 3794
rect 1028 3754 1038 3794
rect 978 3694 1038 3754
rect 978 3654 988 3694
rect 1028 3654 1038 3694
rect 690 3554 700 3594
rect 740 3554 750 3594
rect 832 3626 896 3632
rect 832 3574 838 3626
rect 890 3574 896 3626
rect 832 3568 844 3574
rect 690 3494 750 3554
rect 690 3454 700 3494
rect 740 3454 750 3494
rect 690 3438 750 3454
rect 834 3554 844 3568
rect 884 3568 896 3574
rect 978 3594 1038 3654
rect 884 3554 894 3568
rect 834 3494 894 3554
rect 834 3454 844 3494
rect 884 3454 894 3494
rect 834 3438 894 3454
rect 978 3554 988 3594
rect 1028 3554 1038 3594
rect 978 3494 1038 3554
rect 978 3454 988 3494
rect 1028 3454 1038 3494
rect 978 3438 1038 3454
rect 1266 3794 1326 4000
rect 1266 3754 1276 3794
rect 1316 3754 1326 3794
rect 1266 3694 1326 3754
rect 1266 3654 1276 3694
rect 1316 3654 1326 3694
rect 1266 3594 1326 3654
rect 1410 3794 1470 3844
rect 1410 3754 1420 3794
rect 1460 3754 1470 3794
rect 1410 3694 1470 3754
rect 1410 3654 1420 3694
rect 1460 3654 1470 3694
rect 1410 3632 1470 3654
rect 1554 3794 1614 4000
rect 1554 3754 1564 3794
rect 1604 3754 1614 3794
rect 1554 3694 1614 3754
rect 1554 3654 1564 3694
rect 1604 3654 1614 3694
rect 1266 3554 1276 3594
rect 1316 3554 1326 3594
rect 1408 3626 1472 3632
rect 1408 3574 1414 3626
rect 1466 3574 1472 3626
rect 1408 3568 1420 3574
rect 1266 3494 1326 3554
rect 1266 3454 1276 3494
rect 1316 3454 1326 3494
rect 1266 3438 1326 3454
rect 1410 3554 1420 3568
rect 1460 3568 1472 3574
rect 1554 3594 1614 3654
rect 1460 3554 1470 3568
rect 1410 3494 1470 3554
rect 1410 3454 1420 3494
rect 1460 3454 1470 3494
rect 1410 3438 1470 3454
rect 1554 3554 1564 3594
rect 1604 3554 1614 3594
rect 1554 3494 1614 3554
rect 1554 3454 1564 3494
rect 1604 3454 1614 3494
rect 1554 3438 1614 3454
rect 1842 3794 1902 4000
rect 1842 3754 1852 3794
rect 1892 3754 1902 3794
rect 1842 3694 1902 3754
rect 1842 3654 1852 3694
rect 1892 3654 1902 3694
rect 1842 3594 1902 3654
rect 1986 3794 2046 3844
rect 1986 3754 1996 3794
rect 2036 3754 2046 3794
rect 1986 3694 2046 3754
rect 1986 3654 1996 3694
rect 2036 3654 2046 3694
rect 1986 3632 2046 3654
rect 2130 3794 2190 4000
rect 2130 3754 2140 3794
rect 2180 3754 2190 3794
rect 2130 3694 2190 3754
rect 2130 3654 2140 3694
rect 2180 3654 2190 3694
rect 1842 3554 1852 3594
rect 1892 3554 1902 3594
rect 1984 3626 2048 3632
rect 1984 3574 1990 3626
rect 2042 3574 2048 3626
rect 1984 3568 1996 3574
rect 1842 3494 1902 3554
rect 1842 3454 1852 3494
rect 1892 3454 1902 3494
rect 1842 3438 1902 3454
rect 1986 3554 1996 3568
rect 2036 3568 2048 3574
rect 2130 3594 2190 3654
rect 2036 3554 2046 3568
rect 1986 3494 2046 3554
rect 1986 3454 1996 3494
rect 2036 3454 2046 3494
rect 1986 3438 2046 3454
rect 2130 3554 2140 3594
rect 2180 3554 2190 3594
rect 2130 3494 2190 3554
rect 2130 3454 2140 3494
rect 2180 3454 2190 3494
rect 2130 3438 2190 3454
rect 2418 3794 2478 4000
rect 2418 3754 2428 3794
rect 2468 3754 2478 3794
rect 2418 3694 2478 3754
rect 2418 3654 2428 3694
rect 2468 3654 2478 3694
rect 2418 3594 2478 3654
rect 2562 3794 2622 3844
rect 2562 3754 2572 3794
rect 2612 3754 2622 3794
rect 2562 3694 2622 3754
rect 2562 3654 2572 3694
rect 2612 3654 2622 3694
rect 2562 3632 2622 3654
rect 2706 3794 2766 4000
rect 2706 3754 2716 3794
rect 2756 3754 2766 3794
rect 2706 3694 2766 3754
rect 2706 3654 2716 3694
rect 2756 3654 2766 3694
rect 2418 3554 2428 3594
rect 2468 3554 2478 3594
rect 2560 3626 2624 3632
rect 2560 3574 2566 3626
rect 2618 3574 2624 3626
rect 2560 3568 2572 3574
rect 2418 3494 2478 3554
rect 2418 3454 2428 3494
rect 2468 3454 2478 3494
rect 2418 3438 2478 3454
rect 2562 3554 2572 3568
rect 2612 3568 2624 3574
rect 2706 3594 2766 3654
rect 2612 3554 2622 3568
rect 2562 3494 2622 3554
rect 2562 3454 2572 3494
rect 2612 3454 2622 3494
rect 2562 3438 2622 3454
rect 2706 3554 2716 3594
rect 2756 3554 2766 3594
rect 2706 3494 2766 3554
rect 2706 3454 2716 3494
rect 2756 3454 2766 3494
rect 2706 3438 2766 3454
rect 2994 3794 3054 4000
rect 2994 3754 3004 3794
rect 3044 3754 3054 3794
rect 2994 3694 3054 3754
rect 2994 3654 3004 3694
rect 3044 3654 3054 3694
rect 2994 3594 3054 3654
rect 3138 3794 3198 3844
rect 3138 3754 3148 3794
rect 3188 3754 3198 3794
rect 3138 3694 3198 3754
rect 3138 3654 3148 3694
rect 3188 3654 3198 3694
rect 3138 3632 3198 3654
rect 3282 3794 3342 4000
rect 3282 3754 3292 3794
rect 3332 3754 3342 3794
rect 3282 3694 3342 3754
rect 3282 3654 3292 3694
rect 3332 3654 3342 3694
rect 2994 3554 3004 3594
rect 3044 3554 3054 3594
rect 3136 3626 3200 3632
rect 3136 3574 3142 3626
rect 3194 3574 3200 3626
rect 3136 3568 3148 3574
rect 2994 3494 3054 3554
rect 2994 3454 3004 3494
rect 3044 3454 3054 3494
rect 2994 3438 3054 3454
rect 3138 3554 3148 3568
rect 3188 3568 3200 3574
rect 3282 3594 3342 3654
rect 3188 3554 3198 3568
rect 3138 3494 3198 3554
rect 3138 3454 3148 3494
rect 3188 3454 3198 3494
rect 3138 3438 3198 3454
rect 3282 3554 3292 3594
rect 3332 3554 3342 3594
rect 3282 3494 3342 3554
rect 3570 3704 3630 4000
rect 3570 3552 3580 3704
rect 3620 3552 3630 3704
rect 3714 3704 3774 3844
rect 3714 3632 3724 3704
rect 3712 3626 3724 3632
rect 3764 3632 3774 3704
rect 3858 3704 3918 4000
rect 3764 3626 3776 3632
rect 3712 3574 3718 3626
rect 3770 3574 3776 3626
rect 3712 3568 3724 3574
rect 3570 3528 3630 3552
rect 3714 3552 3724 3568
rect 3764 3568 3776 3574
rect 3764 3552 3774 3568
rect 3714 3528 3774 3552
rect 3858 3552 3868 3704
rect 3908 3552 3918 3704
rect 3858 3528 3918 3552
rect 4146 3794 4206 4000
rect 4146 3754 4156 3794
rect 4196 3754 4206 3794
rect 4146 3694 4206 3754
rect 4146 3654 4156 3694
rect 4196 3654 4206 3694
rect 4146 3594 4206 3654
rect 4290 3794 4350 3844
rect 4290 3754 4300 3794
rect 4340 3754 4350 3794
rect 4290 3694 4350 3754
rect 4290 3654 4300 3694
rect 4340 3654 4350 3694
rect 4290 3632 4350 3654
rect 4434 3794 4494 4000
rect 4434 3754 4444 3794
rect 4484 3754 4494 3794
rect 4434 3694 4494 3754
rect 4434 3654 4444 3694
rect 4484 3654 4494 3694
rect 4146 3554 4156 3594
rect 4196 3554 4206 3594
rect 4288 3626 4352 3632
rect 4288 3574 4294 3626
rect 4346 3574 4352 3626
rect 4288 3568 4300 3574
rect 3282 3454 3292 3494
rect 3332 3454 3342 3494
rect 3282 3438 3342 3454
rect 4146 3494 4206 3554
rect 4146 3454 4156 3494
rect 4196 3454 4206 3494
rect 4146 3438 4206 3454
rect 4290 3554 4300 3568
rect 4340 3568 4352 3574
rect 4434 3594 4494 3654
rect 4340 3554 4350 3568
rect 4290 3494 4350 3554
rect 4290 3454 4300 3494
rect 4340 3454 4350 3494
rect 4290 3438 4350 3454
rect 4434 3554 4444 3594
rect 4484 3554 4494 3594
rect 4434 3494 4494 3554
rect 4434 3454 4444 3494
rect 4484 3454 4494 3494
rect 4434 3438 4494 3454
rect 4722 3794 4782 4000
rect 4722 3754 4732 3794
rect 4772 3754 4782 3794
rect 4722 3694 4782 3754
rect 4722 3654 4732 3694
rect 4772 3654 4782 3694
rect 4722 3594 4782 3654
rect 4866 3794 4926 3844
rect 4866 3754 4876 3794
rect 4916 3754 4926 3794
rect 4866 3694 4926 3754
rect 4866 3654 4876 3694
rect 4916 3654 4926 3694
rect 4866 3632 4926 3654
rect 5010 3794 5070 4000
rect 5010 3754 5020 3794
rect 5060 3754 5070 3794
rect 5010 3694 5070 3754
rect 5010 3654 5020 3694
rect 5060 3654 5070 3694
rect 4722 3554 4732 3594
rect 4772 3554 4782 3594
rect 4864 3626 4928 3632
rect 4864 3574 4870 3626
rect 4922 3574 4928 3626
rect 4864 3568 4876 3574
rect 4722 3494 4782 3554
rect 4722 3454 4732 3494
rect 4772 3454 4782 3494
rect 4722 3438 4782 3454
rect 4866 3554 4876 3568
rect 4916 3568 4928 3574
rect 5010 3594 5070 3654
rect 4916 3554 4926 3568
rect 4866 3494 4926 3554
rect 4866 3454 4876 3494
rect 4916 3454 4926 3494
rect 4866 3438 4926 3454
rect 5010 3554 5020 3594
rect 5060 3554 5070 3594
rect 5010 3494 5070 3554
rect 5010 3454 5020 3494
rect 5060 3454 5070 3494
rect 5010 3438 5070 3454
rect 5298 3794 5358 4000
rect 5298 3754 5308 3794
rect 5348 3754 5358 3794
rect 5298 3694 5358 3754
rect 5298 3654 5308 3694
rect 5348 3654 5358 3694
rect 5298 3594 5358 3654
rect 5442 3794 5502 3844
rect 5442 3754 5452 3794
rect 5492 3754 5502 3794
rect 5442 3694 5502 3754
rect 5442 3654 5452 3694
rect 5492 3654 5502 3694
rect 5442 3632 5502 3654
rect 5586 3794 5646 4000
rect 5586 3754 5596 3794
rect 5636 3754 5646 3794
rect 5586 3694 5646 3754
rect 5586 3654 5596 3694
rect 5636 3654 5646 3694
rect 5298 3554 5308 3594
rect 5348 3554 5358 3594
rect 5440 3626 5504 3632
rect 5440 3574 5446 3626
rect 5498 3574 5504 3626
rect 5440 3568 5452 3574
rect 5298 3494 5358 3554
rect 5298 3454 5308 3494
rect 5348 3454 5358 3494
rect 5298 3438 5358 3454
rect 5442 3554 5452 3568
rect 5492 3568 5504 3574
rect 5586 3594 5646 3654
rect 5874 3794 5934 3844
rect 5874 3754 5884 3794
rect 5924 3754 5934 3794
rect 6018 3794 6078 3844
rect 6018 3776 6028 3794
rect 5874 3694 5934 3754
rect 6016 3770 6028 3776
rect 6068 3776 6078 3794
rect 6162 3794 6222 3844
rect 6068 3770 6080 3776
rect 6016 3718 6022 3770
rect 6074 3718 6080 3770
rect 6016 3712 6080 3718
rect 6162 3754 6172 3794
rect 6212 3754 6222 3794
rect 5874 3654 5884 3694
rect 5924 3654 5934 3694
rect 5874 3632 5934 3654
rect 6018 3694 6078 3712
rect 6018 3654 6028 3694
rect 6068 3654 6078 3694
rect 5492 3554 5502 3568
rect 5442 3494 5502 3554
rect 5442 3454 5452 3494
rect 5492 3454 5502 3494
rect 5442 3438 5502 3454
rect 5586 3554 5596 3594
rect 5636 3554 5646 3594
rect 5872 3626 5936 3632
rect 5872 3574 5878 3626
rect 5930 3574 5936 3626
rect 5872 3568 5884 3574
rect 5586 3494 5646 3554
rect 5586 3454 5596 3494
rect 5636 3454 5646 3494
rect 5586 3438 5646 3454
rect 5874 3554 5884 3568
rect 5924 3568 5936 3574
rect 6018 3594 6078 3654
rect 6162 3694 6222 3754
rect 6162 3654 6172 3694
rect 6212 3654 6222 3694
rect 6162 3632 6222 3654
rect 6450 3794 6510 4000
rect 6450 3754 6460 3794
rect 6500 3754 6510 3794
rect 6450 3694 6510 3754
rect 6450 3654 6460 3694
rect 6500 3654 6510 3694
rect 5924 3554 5934 3568
rect 5874 3494 5934 3554
rect 5874 3454 5884 3494
rect 5924 3454 5934 3494
rect 5874 3438 5934 3454
rect 6018 3554 6028 3594
rect 6068 3554 6078 3594
rect 6160 3626 6224 3632
rect 6160 3574 6166 3626
rect 6218 3574 6224 3626
rect 6160 3568 6172 3574
rect 6018 3494 6078 3554
rect 6018 3454 6028 3494
rect 6068 3454 6078 3494
rect 6018 3438 6078 3454
rect 6162 3554 6172 3568
rect 6212 3568 6224 3574
rect 6450 3594 6510 3654
rect 6212 3554 6222 3568
rect 6162 3494 6222 3554
rect 6162 3454 6172 3494
rect 6212 3454 6222 3494
rect 6162 3438 6222 3454
rect 6450 3554 6460 3594
rect 6500 3554 6510 3594
rect 6450 3494 6510 3554
rect 6450 3454 6460 3494
rect 6500 3454 6510 3494
rect 6450 3438 6510 3454
rect 6594 3794 6654 3844
rect 6594 3754 6604 3794
rect 6644 3754 6654 3794
rect 6738 3794 6798 3844
rect 6738 3776 6748 3794
rect 6594 3694 6654 3754
rect 6736 3770 6748 3776
rect 6788 3776 6798 3794
rect 6788 3770 6800 3776
rect 6736 3718 6742 3770
rect 6794 3718 6800 3770
rect 6736 3712 6800 3718
rect 6594 3654 6604 3694
rect 6644 3654 6654 3694
rect 6594 3594 6654 3654
rect 6594 3554 6604 3594
rect 6644 3554 6654 3594
rect 6594 3494 6654 3554
rect 6594 3454 6604 3494
rect 6644 3454 6654 3494
rect 6594 3438 6654 3454
rect 6738 3694 6798 3712
rect 6738 3654 6748 3694
rect 6788 3654 6798 3694
rect 6738 3594 6798 3654
rect 6738 3554 6748 3594
rect 6788 3554 6798 3594
rect 6738 3494 6798 3554
rect 7026 3704 7086 4000
rect 7026 3552 7036 3704
rect 7076 3552 7086 3704
rect 7170 3704 7230 3844
rect 7170 3632 7180 3704
rect 7168 3626 7180 3632
rect 7220 3632 7230 3704
rect 7314 3704 7374 4000
rect 7220 3626 7232 3632
rect 7168 3574 7174 3626
rect 7226 3574 7232 3626
rect 7168 3568 7180 3574
rect 7026 3528 7086 3552
rect 7170 3552 7180 3568
rect 7220 3568 7232 3574
rect 7220 3552 7230 3568
rect 7170 3528 7230 3552
rect 7314 3552 7324 3704
rect 7364 3552 7374 3704
rect 7314 3528 7374 3552
rect 7602 3794 7662 4000
rect 7602 3754 7612 3794
rect 7652 3754 7662 3794
rect 7602 3694 7662 3754
rect 7602 3654 7612 3694
rect 7652 3654 7662 3694
rect 7602 3594 7662 3654
rect 7746 3794 7806 3844
rect 7746 3754 7756 3794
rect 7796 3754 7806 3794
rect 7746 3694 7806 3754
rect 7746 3654 7756 3694
rect 7796 3654 7806 3694
rect 7746 3632 7806 3654
rect 7890 3794 7950 4000
rect 7890 3754 7900 3794
rect 7940 3754 7950 3794
rect 7890 3694 7950 3754
rect 7890 3654 7900 3694
rect 7940 3654 7950 3694
rect 7602 3554 7612 3594
rect 7652 3554 7662 3594
rect 7744 3626 7808 3632
rect 7744 3574 7750 3626
rect 7802 3574 7808 3626
rect 7744 3568 7756 3574
rect 6738 3454 6748 3494
rect 6788 3454 6798 3494
rect 6738 3438 6798 3454
rect 7602 3494 7662 3554
rect 7602 3454 7612 3494
rect 7652 3454 7662 3494
rect 7602 3438 7662 3454
rect 7746 3554 7756 3568
rect 7796 3568 7808 3574
rect 7890 3594 7950 3654
rect 7796 3554 7806 3568
rect 7746 3494 7806 3554
rect 7746 3454 7756 3494
rect 7796 3454 7806 3494
rect 7746 3438 7806 3454
rect 7890 3554 7900 3594
rect 7940 3554 7950 3594
rect 7890 3494 7950 3554
rect 7890 3454 7900 3494
rect 7940 3454 7950 3494
rect 7890 3438 7950 3454
rect 8178 3794 8238 4000
rect 8178 3754 8188 3794
rect 8228 3754 8238 3794
rect 8178 3694 8238 3754
rect 8178 3654 8188 3694
rect 8228 3654 8238 3694
rect 8178 3594 8238 3654
rect 8322 3794 8382 3844
rect 8322 3754 8332 3794
rect 8372 3754 8382 3794
rect 8322 3694 8382 3754
rect 8322 3654 8332 3694
rect 8372 3654 8382 3694
rect 8322 3632 8382 3654
rect 8466 3794 8526 4000
rect 8466 3754 8476 3794
rect 8516 3754 8526 3794
rect 8466 3694 8526 3754
rect 8466 3654 8476 3694
rect 8516 3654 8526 3694
rect 8178 3554 8188 3594
rect 8228 3554 8238 3594
rect 8320 3626 8384 3632
rect 8320 3574 8326 3626
rect 8378 3574 8384 3626
rect 8320 3568 8332 3574
rect 8178 3494 8238 3554
rect 8178 3454 8188 3494
rect 8228 3454 8238 3494
rect 8178 3438 8238 3454
rect 8322 3554 8332 3568
rect 8372 3568 8384 3574
rect 8466 3594 8526 3654
rect 8754 3794 8814 3844
rect 8754 3754 8764 3794
rect 8804 3754 8814 3794
rect 8898 3794 8958 3844
rect 8898 3776 8908 3794
rect 8754 3694 8814 3754
rect 8896 3770 8908 3776
rect 8948 3776 8958 3794
rect 9042 3794 9102 3844
rect 8948 3770 8960 3776
rect 8896 3718 8902 3770
rect 8954 3718 8960 3770
rect 8896 3712 8960 3718
rect 9042 3754 9052 3794
rect 9092 3754 9102 3794
rect 8754 3654 8764 3694
rect 8804 3654 8814 3694
rect 8754 3632 8814 3654
rect 8898 3694 8958 3712
rect 8898 3654 8908 3694
rect 8948 3654 8958 3694
rect 8372 3554 8382 3568
rect 8322 3494 8382 3554
rect 8322 3454 8332 3494
rect 8372 3454 8382 3494
rect 8322 3438 8382 3454
rect 8466 3554 8476 3594
rect 8516 3554 8526 3594
rect 8752 3626 8816 3632
rect 8752 3574 8758 3626
rect 8810 3574 8816 3626
rect 8752 3568 8764 3574
rect 8466 3494 8526 3554
rect 8466 3454 8476 3494
rect 8516 3454 8526 3494
rect 8466 3438 8526 3454
rect 8754 3554 8764 3568
rect 8804 3568 8816 3574
rect 8898 3594 8958 3654
rect 9042 3694 9102 3754
rect 9042 3654 9052 3694
rect 9092 3654 9102 3694
rect 9042 3632 9102 3654
rect 9330 3794 9390 4000
rect 9330 3754 9340 3794
rect 9380 3754 9390 3794
rect 9330 3694 9390 3754
rect 9330 3654 9340 3694
rect 9380 3654 9390 3694
rect 8804 3554 8814 3568
rect 8754 3494 8814 3554
rect 8754 3454 8764 3494
rect 8804 3454 8814 3494
rect 8754 3438 8814 3454
rect 8898 3554 8908 3594
rect 8948 3554 8958 3594
rect 9040 3626 9104 3632
rect 9040 3574 9046 3626
rect 9098 3574 9104 3626
rect 9040 3568 9052 3574
rect 8898 3494 8958 3554
rect 8898 3454 8908 3494
rect 8948 3454 8958 3494
rect 8898 3438 8958 3454
rect 9042 3554 9052 3568
rect 9092 3568 9104 3574
rect 9330 3594 9390 3654
rect 9092 3554 9102 3568
rect 9042 3494 9102 3554
rect 9042 3454 9052 3494
rect 9092 3454 9102 3494
rect 9042 3438 9102 3454
rect 9330 3554 9340 3594
rect 9380 3554 9390 3594
rect 9330 3494 9390 3554
rect 9330 3454 9340 3494
rect 9380 3454 9390 3494
rect 9330 3438 9390 3454
rect 9474 3794 9534 3844
rect 9474 3754 9484 3794
rect 9524 3754 9534 3794
rect 9618 3794 9678 3844
rect 9618 3776 9628 3794
rect 9474 3694 9534 3754
rect 9616 3770 9628 3776
rect 9668 3776 9678 3794
rect 10194 3794 10254 4000
rect 9668 3770 9680 3776
rect 9616 3718 9622 3770
rect 9674 3718 9680 3770
rect 9616 3712 9680 3718
rect 10194 3754 10204 3794
rect 10244 3754 10254 3794
rect 9474 3654 9484 3694
rect 9524 3654 9534 3694
rect 9474 3594 9534 3654
rect 9474 3554 9484 3594
rect 9524 3554 9534 3594
rect 9474 3494 9534 3554
rect 9474 3454 9484 3494
rect 9524 3454 9534 3494
rect 9474 3438 9534 3454
rect 9618 3694 9678 3712
rect 9618 3654 9628 3694
rect 9668 3654 9678 3694
rect 9618 3594 9678 3654
rect 9618 3554 9628 3594
rect 9668 3554 9678 3594
rect 9618 3494 9678 3554
rect 9618 3454 9628 3494
rect 9668 3454 9678 3494
rect 9618 3438 9678 3454
rect 10194 3694 10254 3754
rect 10194 3654 10204 3694
rect 10244 3654 10254 3694
rect 10194 3594 10254 3654
rect 10338 3794 10398 3844
rect 10338 3754 10348 3794
rect 10388 3754 10398 3794
rect 10338 3694 10398 3754
rect 10338 3654 10348 3694
rect 10388 3654 10398 3694
rect 10338 3632 10398 3654
rect 10482 3794 10542 4000
rect 10482 3754 10492 3794
rect 10532 3754 10542 3794
rect 10482 3694 10542 3754
rect 10482 3654 10492 3694
rect 10532 3654 10542 3694
rect 10194 3554 10204 3594
rect 10244 3554 10254 3594
rect 10336 3626 10400 3632
rect 10336 3574 10342 3626
rect 10394 3574 10400 3626
rect 10336 3568 10348 3574
rect 10194 3494 10254 3554
rect 10194 3454 10204 3494
rect 10244 3454 10254 3494
rect 10194 3438 10254 3454
rect 10338 3554 10348 3568
rect 10388 3568 10400 3574
rect 10482 3594 10542 3654
rect 10388 3554 10398 3568
rect 10338 3494 10398 3554
rect 10338 3454 10348 3494
rect 10388 3454 10398 3494
rect 10338 3438 10398 3454
rect 10482 3554 10492 3594
rect 10532 3554 10542 3594
rect 10482 3494 10542 3554
rect 10482 3454 10492 3494
rect 10532 3454 10542 3494
rect 10482 3438 10542 3454
rect 10770 3794 10830 4000
rect 10770 3754 10780 3794
rect 10820 3754 10830 3794
rect 10770 3694 10830 3754
rect 10770 3654 10780 3694
rect 10820 3654 10830 3694
rect 10770 3594 10830 3654
rect 10914 3794 10974 3844
rect 10914 3754 10924 3794
rect 10964 3754 10974 3794
rect 10914 3694 10974 3754
rect 10914 3654 10924 3694
rect 10964 3654 10974 3694
rect 10914 3632 10974 3654
rect 11058 3794 11118 4000
rect 11058 3754 11068 3794
rect 11108 3754 11118 3794
rect 11058 3694 11118 3754
rect 11058 3654 11068 3694
rect 11108 3654 11118 3694
rect 10770 3554 10780 3594
rect 10820 3554 10830 3594
rect 10912 3626 10976 3632
rect 10912 3574 10918 3626
rect 10970 3574 10976 3626
rect 10912 3568 10924 3574
rect 10770 3494 10830 3554
rect 10770 3454 10780 3494
rect 10820 3454 10830 3494
rect 10770 3438 10830 3454
rect 10914 3554 10924 3568
rect 10964 3568 10976 3574
rect 11058 3594 11118 3654
rect 10964 3554 10974 3568
rect 10914 3494 10974 3554
rect 10914 3454 10924 3494
rect 10964 3454 10974 3494
rect 10914 3438 10974 3454
rect 11058 3554 11068 3594
rect 11108 3554 11118 3594
rect 11058 3494 11118 3554
rect 11346 3704 11406 4000
rect 11346 3552 11356 3704
rect 11396 3552 11406 3704
rect 11490 3704 11550 3844
rect 11490 3632 11500 3704
rect 11488 3626 11500 3632
rect 11540 3632 11550 3704
rect 11634 3704 11694 4000
rect 11540 3626 11552 3632
rect 11488 3574 11494 3626
rect 11546 3574 11552 3626
rect 11488 3568 11500 3574
rect 11346 3528 11406 3552
rect 11490 3552 11500 3568
rect 11540 3568 11552 3574
rect 11540 3552 11550 3568
rect 11490 3528 11550 3552
rect 11634 3552 11644 3704
rect 11684 3552 11694 3704
rect 11634 3528 11694 3552
rect 11922 3794 11982 4000
rect 11922 3754 11932 3794
rect 11972 3754 11982 3794
rect 11922 3694 11982 3754
rect 11922 3654 11932 3694
rect 11972 3654 11982 3694
rect 11922 3594 11982 3654
rect 12066 3794 12126 3844
rect 12066 3754 12076 3794
rect 12116 3754 12126 3794
rect 12066 3694 12126 3754
rect 12066 3654 12076 3694
rect 12116 3654 12126 3694
rect 12066 3632 12126 3654
rect 12210 3794 12270 4000
rect 12210 3754 12220 3794
rect 12260 3754 12270 3794
rect 12498 3794 12558 3844
rect 12498 3776 12508 3794
rect 12210 3694 12270 3754
rect 12496 3770 12508 3776
rect 12548 3776 12558 3794
rect 12642 3794 12702 3844
rect 12548 3770 12560 3776
rect 12496 3718 12502 3770
rect 12554 3718 12560 3770
rect 12496 3712 12560 3718
rect 12642 3754 12652 3794
rect 12692 3754 12702 3794
rect 12786 3794 12846 3844
rect 12786 3776 12796 3794
rect 12210 3654 12220 3694
rect 12260 3654 12270 3694
rect 11922 3554 11932 3594
rect 11972 3554 11982 3594
rect 12064 3626 12128 3632
rect 12064 3574 12070 3626
rect 12122 3574 12128 3626
rect 12064 3568 12076 3574
rect 11058 3454 11068 3494
rect 11108 3454 11118 3494
rect 11058 3438 11118 3454
rect 11922 3494 11982 3554
rect 11922 3454 11932 3494
rect 11972 3454 11982 3494
rect 11922 3438 11982 3454
rect 12066 3554 12076 3568
rect 12116 3568 12128 3574
rect 12210 3594 12270 3654
rect 12116 3554 12126 3568
rect 12066 3494 12126 3554
rect 12066 3454 12076 3494
rect 12116 3454 12126 3494
rect 12066 3438 12126 3454
rect 12210 3554 12220 3594
rect 12260 3554 12270 3594
rect 12210 3494 12270 3554
rect 12210 3454 12220 3494
rect 12260 3454 12270 3494
rect 12210 3438 12270 3454
rect 12498 3694 12558 3712
rect 12498 3654 12508 3694
rect 12548 3654 12558 3694
rect 12498 3594 12558 3654
rect 12642 3694 12702 3754
rect 12784 3770 12796 3776
rect 12836 3776 12846 3794
rect 13650 3794 13710 3844
rect 13650 3776 13660 3794
rect 12836 3770 12848 3776
rect 12784 3718 12790 3770
rect 12842 3718 12848 3770
rect 12784 3712 12848 3718
rect 13648 3770 13660 3776
rect 13700 3776 13710 3794
rect 13794 3794 13854 3844
rect 13700 3770 13712 3776
rect 13648 3718 13654 3770
rect 13706 3718 13712 3770
rect 13648 3712 13712 3718
rect 13794 3754 13804 3794
rect 13844 3754 13854 3794
rect 13938 3794 13998 3844
rect 13938 3776 13948 3794
rect 12642 3654 12652 3694
rect 12692 3654 12702 3694
rect 12642 3632 12702 3654
rect 12786 3694 12846 3712
rect 12786 3654 12796 3694
rect 12836 3654 12846 3694
rect 12498 3554 12508 3594
rect 12548 3554 12558 3594
rect 12640 3626 12704 3632
rect 12640 3574 12646 3626
rect 12698 3574 12704 3626
rect 12640 3568 12652 3574
rect 12498 3494 12558 3554
rect 12498 3454 12508 3494
rect 12548 3454 12558 3494
rect 12498 3438 12558 3454
rect 12642 3554 12652 3568
rect 12692 3568 12704 3574
rect 12786 3594 12846 3654
rect 12692 3554 12702 3568
rect 12642 3494 12702 3554
rect 12642 3454 12652 3494
rect 12692 3454 12702 3494
rect 12642 3438 12702 3454
rect 12786 3554 12796 3594
rect 12836 3554 12846 3594
rect 12786 3494 12846 3554
rect 12786 3454 12796 3494
rect 12836 3454 12846 3494
rect 12786 3438 12846 3454
rect 13650 3694 13710 3712
rect 13650 3654 13660 3694
rect 13700 3654 13710 3694
rect 13650 3594 13710 3654
rect 13794 3694 13854 3754
rect 13936 3770 13948 3776
rect 13988 3776 13998 3794
rect 14226 3794 14286 4000
rect 13988 3770 14000 3776
rect 13936 3718 13942 3770
rect 13994 3718 14000 3770
rect 13936 3712 14000 3718
rect 14226 3754 14236 3794
rect 14276 3754 14286 3794
rect 13794 3654 13804 3694
rect 13844 3654 13854 3694
rect 13794 3632 13854 3654
rect 13938 3694 13998 3712
rect 13938 3654 13948 3694
rect 13988 3654 13998 3694
rect 13650 3554 13660 3594
rect 13700 3554 13710 3594
rect 13792 3626 13856 3632
rect 13792 3574 13798 3626
rect 13850 3574 13856 3626
rect 13792 3568 13804 3574
rect 13650 3494 13710 3554
rect 13650 3454 13660 3494
rect 13700 3454 13710 3494
rect 13650 3438 13710 3454
rect 13794 3554 13804 3568
rect 13844 3568 13856 3574
rect 13938 3594 13998 3654
rect 13844 3554 13854 3568
rect 13794 3494 13854 3554
rect 13794 3454 13804 3494
rect 13844 3454 13854 3494
rect 13794 3438 13854 3454
rect 13938 3554 13948 3594
rect 13988 3554 13998 3594
rect 13938 3494 13998 3554
rect 13938 3454 13948 3494
rect 13988 3454 13998 3494
rect 13938 3438 13998 3454
rect 14226 3694 14286 3754
rect 14226 3654 14236 3694
rect 14276 3654 14286 3694
rect 14226 3594 14286 3654
rect 14370 3794 14430 3844
rect 14370 3754 14380 3794
rect 14420 3754 14430 3794
rect 14370 3694 14430 3754
rect 14370 3654 14380 3694
rect 14420 3654 14430 3694
rect 14370 3632 14430 3654
rect 14514 3794 14574 4000
rect 14514 3754 14524 3794
rect 14564 3754 14574 3794
rect 14514 3694 14574 3754
rect 14514 3654 14524 3694
rect 14564 3654 14574 3694
rect 14226 3554 14236 3594
rect 14276 3554 14286 3594
rect 14368 3626 14432 3632
rect 14368 3574 14374 3626
rect 14426 3574 14432 3626
rect 14368 3568 14380 3574
rect 14226 3494 14286 3554
rect 14226 3454 14236 3494
rect 14276 3454 14286 3494
rect 14226 3438 14286 3454
rect 14370 3554 14380 3568
rect 14420 3568 14432 3574
rect 14514 3594 14574 3654
rect 14420 3554 14430 3568
rect 14370 3494 14430 3554
rect 14370 3454 14380 3494
rect 14420 3454 14430 3494
rect 14370 3438 14430 3454
rect 14514 3554 14524 3594
rect 14564 3554 14574 3594
rect 14514 3494 14574 3554
rect 14514 3454 14524 3494
rect 14564 3454 14574 3494
rect 14514 3438 14574 3454
rect 14802 3794 14862 4000
rect 14802 3754 14812 3794
rect 14852 3754 14862 3794
rect 14802 3694 14862 3754
rect 14802 3654 14812 3694
rect 14852 3654 14862 3694
rect 14802 3594 14862 3654
rect 14946 3794 15006 3844
rect 14946 3754 14956 3794
rect 14996 3754 15006 3794
rect 14946 3694 15006 3754
rect 14946 3654 14956 3694
rect 14996 3654 15006 3694
rect 14946 3632 15006 3654
rect 15090 3794 15150 4000
rect 15090 3754 15100 3794
rect 15140 3754 15150 3794
rect 15090 3694 15150 3754
rect 15090 3654 15100 3694
rect 15140 3654 15150 3694
rect 14802 3554 14812 3594
rect 14852 3554 14862 3594
rect 14944 3626 15008 3632
rect 14944 3574 14950 3626
rect 15002 3574 15008 3626
rect 14944 3568 14956 3574
rect 14802 3494 14862 3554
rect 14802 3454 14812 3494
rect 14852 3454 14862 3494
rect 14802 3438 14862 3454
rect 14946 3554 14956 3568
rect 14996 3568 15008 3574
rect 15090 3594 15150 3654
rect 14996 3554 15006 3568
rect 14946 3494 15006 3554
rect 14946 3454 14956 3494
rect 14996 3454 15006 3494
rect 14946 3438 15006 3454
rect 15090 3554 15100 3594
rect 15140 3554 15150 3594
rect 15090 3494 15150 3554
rect 15378 3704 15438 4000
rect 15378 3552 15388 3704
rect 15428 3552 15438 3704
rect 15522 3704 15582 3844
rect 15522 3632 15532 3704
rect 15520 3626 15532 3632
rect 15572 3632 15582 3704
rect 15666 3704 15726 4000
rect 15572 3626 15584 3632
rect 15520 3574 15526 3626
rect 15578 3574 15584 3626
rect 15520 3568 15532 3574
rect 15378 3528 15438 3552
rect 15522 3552 15532 3568
rect 15572 3568 15584 3574
rect 15572 3552 15582 3568
rect 15522 3528 15582 3552
rect 15666 3552 15676 3704
rect 15716 3552 15726 3704
rect 15666 3528 15726 3552
rect 15954 3704 16014 4000
rect 15954 3552 15964 3704
rect 16004 3552 16014 3704
rect 16098 3704 16158 3844
rect 16098 3632 16108 3704
rect 16096 3626 16108 3632
rect 16148 3632 16158 3704
rect 16242 3704 16302 4000
rect 16148 3626 16160 3632
rect 16096 3574 16102 3626
rect 16154 3574 16160 3626
rect 16096 3568 16108 3574
rect 15954 3528 16014 3552
rect 16098 3552 16108 3568
rect 16148 3568 16160 3574
rect 16148 3552 16158 3568
rect 16098 3528 16158 3552
rect 16242 3552 16252 3704
rect 16292 3552 16302 3704
rect 16242 3528 16302 3552
rect 16530 3794 16590 4000
rect 16530 3754 16540 3794
rect 16580 3754 16590 3794
rect 16530 3694 16590 3754
rect 16530 3654 16540 3694
rect 16580 3654 16590 3694
rect 16530 3594 16590 3654
rect 16674 3794 16734 3844
rect 16674 3754 16684 3794
rect 16724 3754 16734 3794
rect 16674 3694 16734 3754
rect 16674 3654 16684 3694
rect 16724 3654 16734 3694
rect 16674 3632 16734 3654
rect 16818 3794 16878 4000
rect 16818 3754 16828 3794
rect 16868 3754 16878 3794
rect 16818 3694 16878 3754
rect 16818 3654 16828 3694
rect 16868 3654 16878 3694
rect 16530 3554 16540 3594
rect 16580 3554 16590 3594
rect 16672 3626 16736 3632
rect 16672 3574 16678 3626
rect 16730 3574 16736 3626
rect 16672 3568 16684 3574
rect 15090 3454 15100 3494
rect 15140 3454 15150 3494
rect 15090 3438 15150 3454
rect 16530 3494 16590 3554
rect 16530 3454 16540 3494
rect 16580 3454 16590 3494
rect 16530 3438 16590 3454
rect 16674 3554 16684 3568
rect 16724 3568 16736 3574
rect 16818 3594 16878 3654
rect 16962 3794 17022 3844
rect 16962 3754 16972 3794
rect 17012 3754 17022 3794
rect 16962 3694 17022 3754
rect 16962 3654 16972 3694
rect 17012 3654 17022 3694
rect 16962 3632 17022 3654
rect 17106 3794 17166 4000
rect 17106 3754 17116 3794
rect 17156 3754 17166 3794
rect 17106 3694 17166 3754
rect 17106 3654 17116 3694
rect 17156 3654 17166 3694
rect 16724 3554 16734 3568
rect 16674 3494 16734 3554
rect 16674 3454 16684 3494
rect 16724 3454 16734 3494
rect 16674 3438 16734 3454
rect 16818 3554 16828 3594
rect 16868 3554 16878 3594
rect 16960 3626 17024 3632
rect 16960 3574 16966 3626
rect 17018 3574 17024 3626
rect 16960 3568 16972 3574
rect 16818 3494 16878 3554
rect 16818 3454 16828 3494
rect 16868 3454 16878 3494
rect 16818 3438 16878 3454
rect 16962 3554 16972 3568
rect 17012 3568 17024 3574
rect 17106 3594 17166 3654
rect 17250 3794 17310 3844
rect 17250 3754 17260 3794
rect 17300 3754 17310 3794
rect 17250 3694 17310 3754
rect 17250 3654 17260 3694
rect 17300 3654 17310 3694
rect 17250 3632 17310 3654
rect 17394 3794 17454 4000
rect 17394 3754 17404 3794
rect 17444 3754 17454 3794
rect 17394 3694 17454 3754
rect 17394 3654 17404 3694
rect 17444 3654 17454 3694
rect 17012 3554 17022 3568
rect 16962 3494 17022 3554
rect 16962 3454 16972 3494
rect 17012 3454 17022 3494
rect 16962 3438 17022 3454
rect 17106 3554 17116 3594
rect 17156 3554 17166 3594
rect 17248 3626 17312 3632
rect 17248 3574 17254 3626
rect 17306 3574 17312 3626
rect 17248 3568 17260 3574
rect 17106 3494 17166 3554
rect 17106 3454 17116 3494
rect 17156 3454 17166 3494
rect 17106 3438 17166 3454
rect 17250 3554 17260 3568
rect 17300 3568 17312 3574
rect 17394 3594 17454 3654
rect 17538 3794 17598 3844
rect 17538 3754 17548 3794
rect 17588 3754 17598 3794
rect 17538 3694 17598 3754
rect 17538 3654 17548 3694
rect 17588 3654 17598 3694
rect 17538 3632 17598 3654
rect 17682 3794 17742 4000
rect 17682 3754 17692 3794
rect 17732 3754 17742 3794
rect 17682 3694 17742 3754
rect 17682 3654 17692 3694
rect 17732 3654 17742 3694
rect 17300 3554 17310 3568
rect 17250 3494 17310 3554
rect 17250 3454 17260 3494
rect 17300 3454 17310 3494
rect 17250 3438 17310 3454
rect 17394 3554 17404 3594
rect 17444 3554 17454 3594
rect 17536 3626 17600 3632
rect 17536 3574 17542 3626
rect 17594 3574 17600 3626
rect 17536 3568 17548 3574
rect 17394 3494 17454 3554
rect 17394 3454 17404 3494
rect 17444 3454 17454 3494
rect 17394 3438 17454 3454
rect 17538 3554 17548 3568
rect 17588 3568 17600 3574
rect 17682 3594 17742 3654
rect 17826 3794 17886 3844
rect 17826 3754 17836 3794
rect 17876 3754 17886 3794
rect 17826 3694 17886 3754
rect 17826 3654 17836 3694
rect 17876 3654 17886 3694
rect 17826 3632 17886 3654
rect 17970 3794 18030 4000
rect 17970 3754 17980 3794
rect 18020 3754 18030 3794
rect 17970 3694 18030 3754
rect 17970 3654 17980 3694
rect 18020 3654 18030 3694
rect 17588 3554 17598 3568
rect 17538 3494 17598 3554
rect 17538 3454 17548 3494
rect 17588 3454 17598 3494
rect 17538 3438 17598 3454
rect 17682 3554 17692 3594
rect 17732 3554 17742 3594
rect 17824 3626 17888 3632
rect 17824 3574 17830 3626
rect 17882 3574 17888 3626
rect 17824 3568 17836 3574
rect 17682 3494 17742 3554
rect 17682 3454 17692 3494
rect 17732 3454 17742 3494
rect 17682 3438 17742 3454
rect 17826 3554 17836 3568
rect 17876 3568 17888 3574
rect 17970 3594 18030 3654
rect 18114 3794 18174 3844
rect 18114 3754 18124 3794
rect 18164 3754 18174 3794
rect 18114 3694 18174 3754
rect 18114 3654 18124 3694
rect 18164 3654 18174 3694
rect 18114 3632 18174 3654
rect 18258 3794 18318 4000
rect 18258 3754 18268 3794
rect 18308 3754 18318 3794
rect 18258 3694 18318 3754
rect 18258 3654 18268 3694
rect 18308 3654 18318 3694
rect 17876 3554 17886 3568
rect 17826 3494 17886 3554
rect 17826 3454 17836 3494
rect 17876 3454 17886 3494
rect 17826 3438 17886 3454
rect 17970 3554 17980 3594
rect 18020 3554 18030 3594
rect 18112 3626 18176 3632
rect 18112 3574 18118 3626
rect 18170 3574 18176 3626
rect 18112 3568 18124 3574
rect 17970 3494 18030 3554
rect 17970 3454 17980 3494
rect 18020 3454 18030 3494
rect 17970 3438 18030 3454
rect 18114 3554 18124 3568
rect 18164 3568 18176 3574
rect 18258 3594 18318 3654
rect 18402 3794 18462 3844
rect 18402 3754 18412 3794
rect 18452 3754 18462 3794
rect 18402 3694 18462 3754
rect 18402 3654 18412 3694
rect 18452 3654 18462 3694
rect 18402 3632 18462 3654
rect 18546 3794 18606 4000
rect 18546 3754 18556 3794
rect 18596 3754 18606 3794
rect 18546 3694 18606 3754
rect 18546 3654 18556 3694
rect 18596 3654 18606 3694
rect 18164 3554 18174 3568
rect 18114 3494 18174 3554
rect 18114 3454 18124 3494
rect 18164 3454 18174 3494
rect 18114 3438 18174 3454
rect 18258 3554 18268 3594
rect 18308 3554 18318 3594
rect 18400 3626 18464 3632
rect 18400 3574 18406 3626
rect 18458 3574 18464 3626
rect 18400 3568 18412 3574
rect 18258 3494 18318 3554
rect 18258 3454 18268 3494
rect 18308 3454 18318 3494
rect 18258 3438 18318 3454
rect 18402 3554 18412 3568
rect 18452 3568 18464 3574
rect 18546 3594 18606 3654
rect 18690 3794 18750 3844
rect 18690 3754 18700 3794
rect 18740 3754 18750 3794
rect 18690 3694 18750 3754
rect 18690 3654 18700 3694
rect 18740 3654 18750 3694
rect 18690 3632 18750 3654
rect 18834 3794 18894 4000
rect 18834 3754 18844 3794
rect 18884 3754 18894 3794
rect 18834 3694 18894 3754
rect 18834 3654 18844 3694
rect 18884 3654 18894 3694
rect 18452 3554 18462 3568
rect 18402 3494 18462 3554
rect 18402 3454 18412 3494
rect 18452 3454 18462 3494
rect 18402 3438 18462 3454
rect 18546 3554 18556 3594
rect 18596 3554 18606 3594
rect 18688 3626 18752 3632
rect 18688 3574 18694 3626
rect 18746 3574 18752 3626
rect 18688 3568 18700 3574
rect 18546 3494 18606 3554
rect 18546 3454 18556 3494
rect 18596 3454 18606 3494
rect 18546 3438 18606 3454
rect 18690 3554 18700 3568
rect 18740 3568 18752 3574
rect 18834 3594 18894 3654
rect 18978 3794 19038 3844
rect 18978 3754 18988 3794
rect 19028 3754 19038 3794
rect 18978 3694 19038 3754
rect 18978 3654 18988 3694
rect 19028 3654 19038 3694
rect 18978 3632 19038 3654
rect 19122 3794 19182 4000
rect 19122 3754 19132 3794
rect 19172 3754 19182 3794
rect 19122 3694 19182 3754
rect 19122 3654 19132 3694
rect 19172 3654 19182 3694
rect 18740 3554 18750 3568
rect 18690 3494 18750 3554
rect 18690 3454 18700 3494
rect 18740 3454 18750 3494
rect 18690 3438 18750 3454
rect 18834 3554 18844 3594
rect 18884 3554 18894 3594
rect 18976 3626 19040 3632
rect 18976 3574 18982 3626
rect 19034 3574 19040 3626
rect 18976 3568 18988 3574
rect 18834 3494 18894 3554
rect 18834 3454 18844 3494
rect 18884 3454 18894 3494
rect 18834 3438 18894 3454
rect 18978 3554 18988 3568
rect 19028 3568 19040 3574
rect 19122 3594 19182 3654
rect 19266 3794 19326 3844
rect 19266 3754 19276 3794
rect 19316 3754 19326 3794
rect 19266 3694 19326 3754
rect 19266 3654 19276 3694
rect 19316 3654 19326 3694
rect 19266 3632 19326 3654
rect 19410 3794 19470 4000
rect 19410 3754 19420 3794
rect 19460 3754 19470 3794
rect 19410 3694 19470 3754
rect 19410 3654 19420 3694
rect 19460 3654 19470 3694
rect 19028 3554 19038 3568
rect 18978 3494 19038 3554
rect 18978 3454 18988 3494
rect 19028 3454 19038 3494
rect 18978 3438 19038 3454
rect 19122 3554 19132 3594
rect 19172 3554 19182 3594
rect 19264 3626 19328 3632
rect 19264 3574 19270 3626
rect 19322 3574 19328 3626
rect 19264 3568 19276 3574
rect 19122 3494 19182 3554
rect 19122 3454 19132 3494
rect 19172 3454 19182 3494
rect 19122 3438 19182 3454
rect 19266 3554 19276 3568
rect 19316 3568 19328 3574
rect 19410 3594 19470 3654
rect 19554 3794 19614 3844
rect 19554 3754 19564 3794
rect 19604 3754 19614 3794
rect 19554 3694 19614 3754
rect 19554 3654 19564 3694
rect 19604 3654 19614 3694
rect 19554 3632 19614 3654
rect 19698 3794 19758 4000
rect 19698 3754 19708 3794
rect 19748 3754 19758 3794
rect 19698 3694 19758 3754
rect 19698 3654 19708 3694
rect 19748 3654 19758 3694
rect 19316 3554 19326 3568
rect 19266 3494 19326 3554
rect 19266 3454 19276 3494
rect 19316 3454 19326 3494
rect 19266 3438 19326 3454
rect 19410 3554 19420 3594
rect 19460 3554 19470 3594
rect 19552 3626 19616 3632
rect 19552 3574 19558 3626
rect 19610 3574 19616 3626
rect 19552 3568 19564 3574
rect 19410 3494 19470 3554
rect 19410 3454 19420 3494
rect 19460 3454 19470 3494
rect 19410 3438 19470 3454
rect 19554 3554 19564 3568
rect 19604 3568 19616 3574
rect 19698 3594 19758 3654
rect 19842 3794 19902 3844
rect 19842 3754 19852 3794
rect 19892 3754 19902 3794
rect 19842 3694 19902 3754
rect 19842 3654 19852 3694
rect 19892 3654 19902 3694
rect 19842 3632 19902 3654
rect 19986 3794 20046 4000
rect 19986 3754 19996 3794
rect 20036 3754 20046 3794
rect 19986 3694 20046 3754
rect 19986 3654 19996 3694
rect 20036 3654 20046 3694
rect 19604 3554 19614 3568
rect 19554 3494 19614 3554
rect 19554 3454 19564 3494
rect 19604 3454 19614 3494
rect 19554 3438 19614 3454
rect 19698 3554 19708 3594
rect 19748 3554 19758 3594
rect 19840 3626 19904 3632
rect 19840 3574 19846 3626
rect 19898 3574 19904 3626
rect 19840 3568 19852 3574
rect 19698 3494 19758 3554
rect 19698 3454 19708 3494
rect 19748 3454 19758 3494
rect 19698 3438 19758 3454
rect 19842 3554 19852 3568
rect 19892 3568 19904 3574
rect 19986 3594 20046 3654
rect 19892 3554 19902 3568
rect 19842 3494 19902 3554
rect 19842 3454 19852 3494
rect 19892 3454 19902 3494
rect 19842 3438 19902 3454
rect 19986 3554 19996 3594
rect 20036 3554 20046 3594
rect 19986 3494 20046 3554
rect 19986 3454 19996 3494
rect 20036 3454 20046 3494
rect 19986 3438 20046 3454
rect 778 3338 952 3348
rect 778 3329 838 3338
rect 778 3295 790 3329
rect 824 3295 838 3329
rect 778 3286 838 3295
rect 890 3329 952 3338
rect 890 3295 898 3329
rect 932 3295 952 3329
rect 890 3286 952 3295
rect 778 3276 952 3286
rect 1354 3338 1528 3348
rect 1354 3329 1414 3338
rect 1354 3295 1366 3329
rect 1400 3295 1414 3329
rect 1354 3286 1414 3295
rect 1466 3329 1528 3338
rect 1466 3295 1474 3329
rect 1508 3295 1528 3329
rect 1466 3286 1528 3295
rect 1354 3276 1528 3286
rect 1930 3338 2104 3348
rect 1930 3329 1990 3338
rect 1930 3295 1942 3329
rect 1976 3295 1990 3329
rect 1930 3286 1990 3295
rect 2042 3329 2104 3338
rect 2042 3295 2050 3329
rect 2084 3295 2104 3329
rect 2042 3286 2104 3295
rect 1930 3276 2104 3286
rect 2506 3338 2680 3348
rect 2506 3329 2566 3338
rect 2506 3295 2518 3329
rect 2552 3295 2566 3329
rect 2506 3286 2566 3295
rect 2618 3329 2680 3338
rect 2618 3295 2626 3329
rect 2660 3295 2680 3329
rect 2618 3286 2680 3295
rect 2506 3276 2680 3286
rect 3080 3338 3254 3348
rect 3080 3329 3142 3338
rect 3080 3295 3100 3329
rect 3134 3295 3142 3329
rect 3080 3286 3142 3295
rect 3194 3329 3254 3338
rect 3194 3295 3208 3329
rect 3242 3295 3254 3329
rect 3194 3286 3254 3295
rect 3080 3276 3254 3286
rect 4232 3338 4406 3348
rect 4232 3329 4294 3338
rect 4232 3295 4252 3329
rect 4286 3295 4294 3329
rect 4232 3286 4294 3295
rect 4346 3329 4406 3338
rect 4346 3295 4360 3329
rect 4394 3295 4406 3329
rect 4346 3286 4406 3295
rect 4232 3276 4406 3286
rect 4808 3338 4982 3348
rect 4808 3329 4870 3338
rect 4808 3295 4828 3329
rect 4862 3295 4870 3329
rect 4808 3286 4870 3295
rect 4922 3329 4982 3338
rect 4922 3295 4936 3329
rect 4970 3295 4982 3329
rect 4922 3286 4982 3295
rect 4808 3276 4982 3286
rect 5384 3338 5558 3348
rect 5384 3329 5446 3338
rect 5384 3295 5404 3329
rect 5438 3295 5446 3329
rect 5384 3286 5446 3295
rect 5498 3329 5558 3338
rect 5498 3295 5512 3329
rect 5546 3295 5558 3329
rect 5498 3286 5558 3295
rect 5384 3276 5558 3286
rect 5960 3338 6134 3348
rect 5960 3329 6022 3338
rect 5960 3295 5980 3329
rect 6014 3295 6022 3329
rect 5960 3286 6022 3295
rect 6074 3329 6134 3338
rect 6074 3295 6088 3329
rect 6122 3295 6134 3329
rect 6074 3286 6134 3295
rect 5960 3276 6134 3286
rect 6446 3330 6536 3348
rect 6446 3294 6468 3330
rect 6504 3294 6536 3330
rect 6446 3276 6536 3294
rect 6710 3338 6800 3348
rect 6710 3286 6742 3338
rect 6794 3286 6800 3338
rect 6710 3276 6800 3286
rect 7688 3338 7862 3348
rect 7688 3329 7750 3338
rect 7688 3295 7708 3329
rect 7742 3295 7750 3329
rect 7688 3286 7750 3295
rect 7802 3329 7862 3338
rect 7802 3295 7816 3329
rect 7850 3295 7862 3329
rect 7802 3286 7862 3295
rect 7688 3276 7862 3286
rect 8264 3338 8438 3348
rect 8264 3329 8326 3338
rect 8264 3295 8284 3329
rect 8318 3295 8326 3329
rect 8264 3286 8326 3295
rect 8378 3329 8438 3338
rect 8378 3295 8392 3329
rect 8426 3295 8438 3329
rect 8378 3286 8438 3295
rect 8264 3276 8438 3286
rect 8840 3338 9014 3348
rect 8840 3329 8902 3338
rect 8840 3295 8860 3329
rect 8894 3295 8902 3329
rect 8840 3286 8902 3295
rect 8954 3329 9014 3338
rect 8954 3295 8968 3329
rect 9002 3295 9014 3329
rect 8954 3286 9014 3295
rect 8840 3276 9014 3286
rect 9326 3330 9416 3348
rect 9326 3294 9348 3330
rect 9384 3294 9416 3330
rect 9326 3276 9416 3294
rect 9590 3338 9680 3348
rect 9590 3286 9622 3338
rect 9674 3286 9680 3338
rect 9590 3276 9680 3286
rect 10280 3338 10454 3348
rect 10280 3329 10342 3338
rect 10280 3295 10300 3329
rect 10334 3295 10342 3329
rect 10280 3286 10342 3295
rect 10394 3329 10454 3338
rect 10394 3295 10408 3329
rect 10442 3295 10454 3329
rect 10394 3286 10454 3295
rect 10280 3276 10454 3286
rect 10856 3338 11030 3348
rect 10856 3329 10918 3338
rect 10856 3295 10876 3329
rect 10910 3295 10918 3329
rect 10856 3286 10918 3295
rect 10970 3329 11030 3338
rect 10970 3295 10984 3329
rect 11018 3295 11030 3329
rect 10970 3286 11030 3295
rect 10856 3276 11030 3286
rect 12008 3338 12182 3348
rect 12008 3329 12070 3338
rect 12008 3295 12028 3329
rect 12062 3295 12070 3329
rect 12008 3286 12070 3295
rect 12122 3329 12182 3338
rect 12122 3295 12136 3329
rect 12170 3295 12182 3329
rect 12122 3286 12182 3295
rect 12008 3276 12182 3286
rect 12584 3338 12758 3348
rect 12584 3329 12646 3338
rect 12584 3295 12604 3329
rect 12638 3295 12646 3329
rect 12584 3286 12646 3295
rect 12698 3329 12758 3338
rect 12698 3295 12712 3329
rect 12746 3295 12758 3329
rect 12698 3286 12758 3295
rect 12584 3276 12758 3286
rect 13736 3338 13910 3348
rect 13736 3329 13798 3338
rect 13736 3295 13756 3329
rect 13790 3295 13798 3329
rect 13736 3286 13798 3295
rect 13850 3329 13910 3338
rect 13850 3295 13864 3329
rect 13898 3295 13910 3329
rect 13850 3286 13910 3295
rect 13736 3276 13910 3286
rect 14312 3338 14486 3348
rect 14312 3329 14374 3338
rect 14312 3295 14332 3329
rect 14366 3295 14374 3329
rect 14312 3286 14374 3295
rect 14426 3329 14486 3338
rect 14426 3295 14440 3329
rect 14474 3295 14486 3329
rect 14426 3286 14486 3295
rect 14312 3276 14486 3286
rect 14888 3338 15062 3348
rect 14888 3329 14950 3338
rect 14888 3295 14908 3329
rect 14942 3295 14950 3329
rect 14888 3286 14950 3295
rect 15002 3329 15062 3338
rect 15002 3295 15016 3329
rect 15050 3295 15062 3329
rect 15002 3286 15062 3295
rect 14888 3276 15062 3286
rect 16618 3338 16792 3348
rect 16618 3329 16678 3338
rect 16618 3295 16630 3329
rect 16664 3295 16678 3329
rect 16618 3286 16678 3295
rect 16730 3329 16792 3338
rect 16730 3295 16738 3329
rect 16772 3295 16792 3329
rect 16730 3286 16792 3295
rect 16618 3276 16792 3286
rect 16906 3338 17080 3348
rect 16906 3329 16966 3338
rect 16906 3295 16918 3329
rect 16952 3295 16966 3329
rect 16906 3286 16966 3295
rect 17018 3329 17080 3338
rect 17018 3295 17026 3329
rect 17060 3295 17080 3329
rect 17018 3286 17080 3295
rect 16906 3276 17080 3286
rect 17194 3338 17368 3348
rect 17194 3329 17254 3338
rect 17194 3295 17206 3329
rect 17240 3295 17254 3329
rect 17194 3286 17254 3295
rect 17306 3329 17368 3338
rect 17306 3295 17314 3329
rect 17348 3295 17368 3329
rect 17306 3286 17368 3295
rect 17194 3276 17368 3286
rect 17482 3338 17656 3348
rect 17482 3329 17542 3338
rect 17482 3295 17494 3329
rect 17528 3295 17542 3329
rect 17482 3286 17542 3295
rect 17594 3329 17656 3338
rect 17594 3295 17602 3329
rect 17636 3295 17656 3329
rect 17594 3286 17656 3295
rect 17482 3276 17656 3286
rect 17770 3338 17944 3348
rect 17770 3329 17830 3338
rect 17770 3295 17782 3329
rect 17816 3295 17830 3329
rect 17770 3286 17830 3295
rect 17882 3329 17944 3338
rect 17882 3295 17890 3329
rect 17924 3295 17944 3329
rect 17882 3286 17944 3295
rect 17770 3276 17944 3286
rect 18058 3338 18232 3348
rect 18058 3329 18118 3338
rect 18058 3295 18070 3329
rect 18104 3295 18118 3329
rect 18058 3286 18118 3295
rect 18170 3329 18232 3338
rect 18170 3295 18178 3329
rect 18212 3295 18232 3329
rect 18170 3286 18232 3295
rect 18058 3276 18232 3286
rect 18346 3338 18520 3348
rect 18346 3329 18406 3338
rect 18346 3295 18358 3329
rect 18392 3295 18406 3329
rect 18346 3286 18406 3295
rect 18458 3329 18520 3338
rect 18458 3295 18466 3329
rect 18500 3295 18520 3329
rect 18458 3286 18520 3295
rect 18346 3276 18520 3286
rect 18634 3338 18808 3348
rect 18634 3329 18694 3338
rect 18634 3295 18646 3329
rect 18680 3295 18694 3329
rect 18634 3286 18694 3295
rect 18746 3329 18808 3338
rect 18746 3295 18754 3329
rect 18788 3295 18808 3329
rect 18746 3286 18808 3295
rect 18634 3276 18808 3286
rect 18922 3338 19096 3348
rect 18922 3329 18982 3338
rect 18922 3295 18934 3329
rect 18968 3295 18982 3329
rect 18922 3286 18982 3295
rect 19034 3329 19096 3338
rect 19034 3295 19042 3329
rect 19076 3295 19096 3329
rect 19034 3286 19096 3295
rect 18922 3276 19096 3286
rect 19210 3338 19384 3348
rect 19210 3329 19270 3338
rect 19210 3295 19222 3329
rect 19256 3295 19270 3329
rect 19210 3286 19270 3295
rect 19322 3329 19384 3338
rect 19322 3295 19330 3329
rect 19364 3295 19384 3329
rect 19322 3286 19384 3295
rect 19210 3276 19384 3286
rect 19498 3338 19672 3348
rect 19498 3329 19558 3338
rect 19498 3295 19510 3329
rect 19544 3295 19558 3329
rect 19498 3286 19558 3295
rect 19610 3329 19672 3338
rect 19610 3295 19618 3329
rect 19652 3295 19672 3329
rect 19610 3286 19672 3295
rect 19498 3276 19672 3286
rect 19786 3338 19960 3348
rect 19786 3329 19846 3338
rect 19786 3295 19798 3329
rect 19832 3295 19846 3329
rect 19786 3286 19846 3295
rect 19898 3329 19960 3338
rect 19898 3295 19906 3329
rect 19940 3295 19960 3329
rect 19898 3286 19960 3295
rect 19786 3276 19960 3286
rect 6450 3056 6510 3276
rect 9330 3056 9390 3276
rect 6448 3050 6512 3056
rect 6448 2998 6454 3050
rect 6506 2998 6512 3050
rect 6448 2992 6512 2998
rect 9328 3050 9392 3056
rect 9328 2998 9334 3050
rect 9386 2998 9392 3050
rect 9328 2992 9392 2998
rect 6450 2772 6510 2992
rect 9330 2772 9390 2992
rect 778 2762 952 2772
rect 778 2753 838 2762
rect 778 2719 790 2753
rect 824 2719 838 2753
rect 778 2710 838 2719
rect 890 2753 952 2762
rect 890 2719 898 2753
rect 932 2719 952 2753
rect 890 2710 952 2719
rect 778 2700 952 2710
rect 1354 2762 1528 2772
rect 1354 2753 1414 2762
rect 1354 2719 1366 2753
rect 1400 2719 1414 2753
rect 1354 2710 1414 2719
rect 1466 2753 1528 2762
rect 1466 2719 1474 2753
rect 1508 2719 1528 2753
rect 1466 2710 1528 2719
rect 1354 2700 1528 2710
rect 1930 2762 2104 2772
rect 1930 2753 1990 2762
rect 1930 2719 1942 2753
rect 1976 2719 1990 2753
rect 1930 2710 1990 2719
rect 2042 2753 2104 2762
rect 2042 2719 2050 2753
rect 2084 2719 2104 2753
rect 2042 2710 2104 2719
rect 1930 2700 2104 2710
rect 2506 2762 2680 2772
rect 2506 2753 2566 2762
rect 2506 2719 2518 2753
rect 2552 2719 2566 2753
rect 2506 2710 2566 2719
rect 2618 2753 2680 2762
rect 2618 2719 2626 2753
rect 2660 2719 2680 2753
rect 2618 2710 2680 2719
rect 2506 2700 2680 2710
rect 3080 2762 3254 2772
rect 3080 2753 3142 2762
rect 3080 2719 3100 2753
rect 3134 2719 3142 2753
rect 3080 2710 3142 2719
rect 3194 2753 3254 2762
rect 3194 2719 3208 2753
rect 3242 2719 3254 2753
rect 3194 2710 3254 2719
rect 3080 2700 3254 2710
rect 4232 2762 4406 2772
rect 4232 2753 4294 2762
rect 4232 2719 4252 2753
rect 4286 2719 4294 2753
rect 4232 2710 4294 2719
rect 4346 2753 4406 2762
rect 4346 2719 4360 2753
rect 4394 2719 4406 2753
rect 4346 2710 4406 2719
rect 4232 2700 4406 2710
rect 4808 2762 4982 2772
rect 4808 2753 4870 2762
rect 4808 2719 4828 2753
rect 4862 2719 4870 2753
rect 4808 2710 4870 2719
rect 4922 2753 4982 2762
rect 4922 2719 4936 2753
rect 4970 2719 4982 2753
rect 4922 2710 4982 2719
rect 4808 2700 4982 2710
rect 5384 2762 5558 2772
rect 5384 2753 5446 2762
rect 5384 2719 5404 2753
rect 5438 2719 5446 2753
rect 5384 2710 5446 2719
rect 5498 2753 5558 2762
rect 5498 2719 5512 2753
rect 5546 2719 5558 2753
rect 5498 2710 5558 2719
rect 5384 2700 5558 2710
rect 5960 2762 6134 2772
rect 5960 2753 6022 2762
rect 5960 2719 5980 2753
rect 6014 2719 6022 2753
rect 5960 2710 6022 2719
rect 6074 2753 6134 2762
rect 6074 2719 6088 2753
rect 6122 2719 6134 2753
rect 6074 2710 6134 2719
rect 5960 2700 6134 2710
rect 6446 2754 6536 2772
rect 6446 2718 6468 2754
rect 6504 2718 6536 2754
rect 6446 2700 6536 2718
rect 6710 2762 6800 2772
rect 6710 2710 6742 2762
rect 6794 2710 6800 2762
rect 6710 2700 6800 2710
rect 7688 2762 7862 2772
rect 7688 2753 7750 2762
rect 7688 2719 7708 2753
rect 7742 2719 7750 2753
rect 7688 2710 7750 2719
rect 7802 2753 7862 2762
rect 7802 2719 7816 2753
rect 7850 2719 7862 2753
rect 7802 2710 7862 2719
rect 7688 2700 7862 2710
rect 8264 2762 8438 2772
rect 8264 2753 8326 2762
rect 8264 2719 8284 2753
rect 8318 2719 8326 2753
rect 8264 2710 8326 2719
rect 8378 2753 8438 2762
rect 8378 2719 8392 2753
rect 8426 2719 8438 2753
rect 8378 2710 8438 2719
rect 8264 2700 8438 2710
rect 8840 2762 9014 2772
rect 8840 2753 8902 2762
rect 8840 2719 8860 2753
rect 8894 2719 8902 2753
rect 8840 2710 8902 2719
rect 8954 2753 9014 2762
rect 8954 2719 8968 2753
rect 9002 2719 9014 2753
rect 8954 2710 9014 2719
rect 8840 2700 9014 2710
rect 9326 2754 9416 2772
rect 9326 2718 9348 2754
rect 9384 2718 9416 2754
rect 9326 2700 9416 2718
rect 9590 2762 9680 2772
rect 9590 2710 9622 2762
rect 9674 2710 9680 2762
rect 9590 2700 9680 2710
rect 10280 2762 10454 2772
rect 10280 2753 10342 2762
rect 10280 2719 10300 2753
rect 10334 2719 10342 2753
rect 10280 2710 10342 2719
rect 10394 2753 10454 2762
rect 10394 2719 10408 2753
rect 10442 2719 10454 2753
rect 10394 2710 10454 2719
rect 10280 2700 10454 2710
rect 10856 2762 11030 2772
rect 10856 2753 10918 2762
rect 10856 2719 10876 2753
rect 10910 2719 10918 2753
rect 10856 2710 10918 2719
rect 10970 2753 11030 2762
rect 10970 2719 10984 2753
rect 11018 2719 11030 2753
rect 10970 2710 11030 2719
rect 10856 2700 11030 2710
rect 12008 2762 12182 2772
rect 12008 2753 12070 2762
rect 12008 2719 12028 2753
rect 12062 2719 12070 2753
rect 12008 2710 12070 2719
rect 12122 2753 12182 2762
rect 12122 2719 12136 2753
rect 12170 2719 12182 2753
rect 12122 2710 12182 2719
rect 12008 2700 12182 2710
rect 12584 2762 12758 2772
rect 12584 2753 12646 2762
rect 12584 2719 12604 2753
rect 12638 2719 12646 2753
rect 12584 2710 12646 2719
rect 12698 2753 12758 2762
rect 12698 2719 12712 2753
rect 12746 2719 12758 2753
rect 12698 2710 12758 2719
rect 12584 2700 12758 2710
rect 13736 2762 13910 2772
rect 13736 2753 13798 2762
rect 13736 2719 13756 2753
rect 13790 2719 13798 2753
rect 13736 2710 13798 2719
rect 13850 2753 13910 2762
rect 13850 2719 13864 2753
rect 13898 2719 13910 2753
rect 13850 2710 13910 2719
rect 13736 2700 13910 2710
rect 14312 2762 14486 2772
rect 14312 2753 14374 2762
rect 14312 2719 14332 2753
rect 14366 2719 14374 2753
rect 14312 2710 14374 2719
rect 14426 2753 14486 2762
rect 14426 2719 14440 2753
rect 14474 2719 14486 2753
rect 14426 2710 14486 2719
rect 14312 2700 14486 2710
rect 14888 2762 15062 2772
rect 14888 2753 14950 2762
rect 14888 2719 14908 2753
rect 14942 2719 14950 2753
rect 14888 2710 14950 2719
rect 15002 2753 15062 2762
rect 15002 2719 15016 2753
rect 15050 2719 15062 2753
rect 15002 2710 15062 2719
rect 14888 2700 15062 2710
rect 16618 2762 16792 2772
rect 16618 2753 16678 2762
rect 16618 2719 16630 2753
rect 16664 2719 16678 2753
rect 16618 2710 16678 2719
rect 16730 2753 16792 2762
rect 16730 2719 16738 2753
rect 16772 2719 16792 2753
rect 16730 2710 16792 2719
rect 16618 2700 16792 2710
rect 16906 2762 17080 2772
rect 16906 2753 16966 2762
rect 16906 2719 16918 2753
rect 16952 2719 16966 2753
rect 16906 2710 16966 2719
rect 17018 2753 17080 2762
rect 17018 2719 17026 2753
rect 17060 2719 17080 2753
rect 17018 2710 17080 2719
rect 16906 2700 17080 2710
rect 17194 2762 17368 2772
rect 17194 2753 17254 2762
rect 17194 2719 17206 2753
rect 17240 2719 17254 2753
rect 17194 2710 17254 2719
rect 17306 2753 17368 2762
rect 17306 2719 17314 2753
rect 17348 2719 17368 2753
rect 17306 2710 17368 2719
rect 17194 2700 17368 2710
rect 17482 2762 17656 2772
rect 17482 2753 17542 2762
rect 17482 2719 17494 2753
rect 17528 2719 17542 2753
rect 17482 2710 17542 2719
rect 17594 2753 17656 2762
rect 17594 2719 17602 2753
rect 17636 2719 17656 2753
rect 17594 2710 17656 2719
rect 17482 2700 17656 2710
rect 17770 2762 17944 2772
rect 17770 2753 17830 2762
rect 17770 2719 17782 2753
rect 17816 2719 17830 2753
rect 17770 2710 17830 2719
rect 17882 2753 17944 2762
rect 17882 2719 17890 2753
rect 17924 2719 17944 2753
rect 17882 2710 17944 2719
rect 17770 2700 17944 2710
rect 18058 2762 18232 2772
rect 18058 2753 18118 2762
rect 18058 2719 18070 2753
rect 18104 2719 18118 2753
rect 18058 2710 18118 2719
rect 18170 2753 18232 2762
rect 18170 2719 18178 2753
rect 18212 2719 18232 2753
rect 18170 2710 18232 2719
rect 18058 2700 18232 2710
rect 18346 2762 18520 2772
rect 18346 2753 18406 2762
rect 18346 2719 18358 2753
rect 18392 2719 18406 2753
rect 18346 2710 18406 2719
rect 18458 2753 18520 2762
rect 18458 2719 18466 2753
rect 18500 2719 18520 2753
rect 18458 2710 18520 2719
rect 18346 2700 18520 2710
rect 18634 2762 18808 2772
rect 18634 2753 18694 2762
rect 18634 2719 18646 2753
rect 18680 2719 18694 2753
rect 18634 2710 18694 2719
rect 18746 2753 18808 2762
rect 18746 2719 18754 2753
rect 18788 2719 18808 2753
rect 18746 2710 18808 2719
rect 18634 2700 18808 2710
rect 18922 2762 19096 2772
rect 18922 2753 18982 2762
rect 18922 2719 18934 2753
rect 18968 2719 18982 2753
rect 18922 2710 18982 2719
rect 19034 2753 19096 2762
rect 19034 2719 19042 2753
rect 19076 2719 19096 2753
rect 19034 2710 19096 2719
rect 18922 2700 19096 2710
rect 19210 2762 19384 2772
rect 19210 2753 19270 2762
rect 19210 2719 19222 2753
rect 19256 2719 19270 2753
rect 19210 2710 19270 2719
rect 19322 2753 19384 2762
rect 19322 2719 19330 2753
rect 19364 2719 19384 2753
rect 19322 2710 19384 2719
rect 19210 2700 19384 2710
rect 19498 2762 19672 2772
rect 19498 2753 19558 2762
rect 19498 2719 19510 2753
rect 19544 2719 19558 2753
rect 19498 2710 19558 2719
rect 19610 2753 19672 2762
rect 19610 2719 19618 2753
rect 19652 2719 19672 2753
rect 19610 2710 19672 2719
rect 19498 2700 19672 2710
rect 19786 2762 19960 2772
rect 19786 2753 19846 2762
rect 19786 2719 19798 2753
rect 19832 2719 19846 2753
rect 19786 2710 19846 2719
rect 19898 2753 19960 2762
rect 19898 2719 19906 2753
rect 19940 2719 19960 2753
rect 19898 2710 19960 2719
rect 19786 2700 19960 2710
rect 114 2588 174 2630
rect 114 2500 124 2588
rect 164 2500 174 2588
rect 114 2048 174 2500
rect 258 2588 318 2630
rect 258 2500 268 2588
rect 308 2500 318 2588
rect 258 2480 318 2500
rect 402 2588 462 2630
rect 402 2500 412 2588
rect 452 2500 462 2588
rect 256 2474 320 2480
rect 256 2422 262 2474
rect 314 2422 320 2474
rect 256 2416 320 2422
rect 258 2302 318 2416
rect 402 2048 462 2500
rect 690 2614 750 2630
rect 690 2574 700 2614
rect 740 2574 750 2614
rect 690 2514 750 2574
rect 690 2474 700 2514
rect 740 2474 750 2514
rect 834 2614 894 2630
rect 834 2574 844 2614
rect 884 2574 894 2614
rect 834 2514 894 2574
rect 834 2480 844 2514
rect 690 2048 750 2474
rect 832 2474 844 2480
rect 884 2480 894 2514
rect 978 2614 1038 2630
rect 978 2574 988 2614
rect 1028 2574 1038 2614
rect 978 2514 1038 2574
rect 884 2474 896 2480
rect 832 2422 838 2474
rect 890 2422 896 2474
rect 832 2416 896 2422
rect 978 2474 988 2514
rect 1028 2474 1038 2514
rect 834 2302 894 2416
rect 978 2048 1038 2474
rect 1266 2614 1326 2630
rect 1266 2574 1276 2614
rect 1316 2574 1326 2614
rect 1266 2514 1326 2574
rect 1266 2474 1276 2514
rect 1316 2474 1326 2514
rect 1410 2614 1470 2630
rect 1410 2574 1420 2614
rect 1460 2574 1470 2614
rect 1410 2514 1470 2574
rect 1410 2480 1420 2514
rect 1266 2048 1326 2474
rect 1408 2474 1420 2480
rect 1460 2480 1470 2514
rect 1554 2614 1614 2630
rect 1554 2574 1564 2614
rect 1604 2574 1614 2614
rect 1554 2514 1614 2574
rect 1460 2474 1472 2480
rect 1408 2422 1414 2474
rect 1466 2422 1472 2474
rect 1408 2416 1472 2422
rect 1554 2474 1564 2514
rect 1604 2474 1614 2514
rect 1410 2302 1470 2416
rect 1554 2048 1614 2474
rect 1842 2614 1902 2630
rect 1842 2574 1852 2614
rect 1892 2574 1902 2614
rect 1842 2514 1902 2574
rect 1842 2474 1852 2514
rect 1892 2474 1902 2514
rect 1986 2614 2046 2630
rect 1986 2574 1996 2614
rect 2036 2574 2046 2614
rect 1986 2514 2046 2574
rect 1986 2480 1996 2514
rect 1842 2048 1902 2474
rect 1984 2474 1996 2480
rect 2036 2480 2046 2514
rect 2130 2614 2190 2630
rect 2130 2574 2140 2614
rect 2180 2574 2190 2614
rect 2130 2514 2190 2574
rect 2036 2474 2048 2480
rect 1984 2422 1990 2474
rect 2042 2422 2048 2474
rect 1984 2416 2048 2422
rect 2130 2474 2140 2514
rect 2180 2474 2190 2514
rect 1986 2302 2046 2416
rect 2130 2048 2190 2474
rect 2418 2614 2478 2630
rect 2418 2574 2428 2614
rect 2468 2574 2478 2614
rect 2418 2514 2478 2574
rect 2418 2474 2428 2514
rect 2468 2474 2478 2514
rect 2562 2614 2622 2630
rect 2562 2574 2572 2614
rect 2612 2574 2622 2614
rect 2562 2514 2622 2574
rect 2562 2480 2572 2514
rect 2418 2048 2478 2474
rect 2560 2474 2572 2480
rect 2612 2480 2622 2514
rect 2706 2614 2766 2630
rect 2706 2574 2716 2614
rect 2756 2574 2766 2614
rect 2706 2514 2766 2574
rect 2612 2474 2624 2480
rect 2560 2422 2566 2474
rect 2618 2422 2624 2474
rect 2560 2416 2624 2422
rect 2706 2474 2716 2514
rect 2756 2474 2766 2514
rect 2562 2302 2622 2416
rect 2706 2048 2766 2474
rect 2994 2614 3054 2630
rect 2994 2574 3004 2614
rect 3044 2574 3054 2614
rect 2994 2514 3054 2574
rect 2994 2474 3004 2514
rect 3044 2474 3054 2514
rect 3138 2614 3198 2630
rect 3138 2574 3148 2614
rect 3188 2574 3198 2614
rect 3138 2514 3198 2574
rect 3138 2480 3148 2514
rect 2994 2048 3054 2474
rect 3136 2474 3148 2480
rect 3188 2480 3198 2514
rect 3282 2614 3342 2630
rect 3282 2574 3292 2614
rect 3332 2574 3342 2614
rect 3282 2514 3342 2574
rect 3188 2474 3200 2480
rect 3136 2422 3142 2474
rect 3194 2422 3200 2474
rect 3136 2416 3200 2422
rect 3282 2474 3292 2514
rect 3332 2474 3342 2514
rect 3138 2302 3198 2416
rect 3282 2048 3342 2474
rect 3570 2588 3630 2630
rect 3570 2500 3580 2588
rect 3620 2500 3630 2588
rect 3570 2048 3630 2500
rect 3714 2588 3774 2630
rect 3714 2500 3724 2588
rect 3764 2500 3774 2588
rect 3714 2480 3774 2500
rect 3858 2588 3918 2630
rect 3858 2500 3868 2588
rect 3908 2500 3918 2588
rect 3712 2474 3776 2480
rect 3712 2422 3718 2474
rect 3770 2422 3776 2474
rect 3712 2416 3776 2422
rect 3714 2302 3774 2416
rect 3858 2048 3918 2500
rect 4146 2614 4206 2630
rect 4146 2574 4156 2614
rect 4196 2574 4206 2614
rect 4146 2514 4206 2574
rect 4146 2474 4156 2514
rect 4196 2474 4206 2514
rect 4290 2614 4350 2630
rect 4290 2574 4300 2614
rect 4340 2574 4350 2614
rect 4290 2514 4350 2574
rect 4290 2480 4300 2514
rect 4146 2048 4206 2474
rect 4288 2474 4300 2480
rect 4340 2480 4350 2514
rect 4434 2614 4494 2630
rect 4434 2574 4444 2614
rect 4484 2574 4494 2614
rect 4434 2514 4494 2574
rect 4340 2474 4352 2480
rect 4288 2422 4294 2474
rect 4346 2422 4352 2474
rect 4288 2416 4352 2422
rect 4434 2474 4444 2514
rect 4484 2474 4494 2514
rect 4290 2302 4350 2416
rect 4434 2048 4494 2474
rect 4722 2614 4782 2630
rect 4722 2574 4732 2614
rect 4772 2574 4782 2614
rect 4722 2514 4782 2574
rect 4722 2474 4732 2514
rect 4772 2474 4782 2514
rect 4866 2614 4926 2630
rect 4866 2574 4876 2614
rect 4916 2574 4926 2614
rect 4866 2514 4926 2574
rect 4866 2480 4876 2514
rect 4722 2048 4782 2474
rect 4864 2474 4876 2480
rect 4916 2480 4926 2514
rect 5010 2614 5070 2630
rect 5010 2574 5020 2614
rect 5060 2574 5070 2614
rect 5010 2514 5070 2574
rect 4916 2474 4928 2480
rect 4864 2422 4870 2474
rect 4922 2422 4928 2474
rect 4864 2416 4928 2422
rect 5010 2474 5020 2514
rect 5060 2474 5070 2514
rect 4866 2302 4926 2416
rect 5010 2048 5070 2474
rect 5298 2614 5358 2630
rect 5298 2574 5308 2614
rect 5348 2574 5358 2614
rect 5298 2514 5358 2574
rect 5298 2474 5308 2514
rect 5348 2474 5358 2514
rect 5442 2614 5502 2630
rect 5442 2574 5452 2614
rect 5492 2574 5502 2614
rect 5442 2514 5502 2574
rect 5442 2480 5452 2514
rect 5298 2048 5358 2474
rect 5440 2474 5452 2480
rect 5492 2480 5502 2514
rect 5586 2614 5646 2630
rect 5586 2574 5596 2614
rect 5636 2574 5646 2614
rect 5586 2514 5646 2574
rect 5492 2474 5504 2480
rect 5440 2422 5446 2474
rect 5498 2422 5504 2474
rect 5440 2416 5504 2422
rect 5586 2474 5596 2514
rect 5636 2474 5646 2514
rect 5874 2614 5934 2630
rect 5874 2574 5884 2614
rect 5924 2574 5934 2614
rect 5874 2514 5934 2574
rect 5874 2480 5884 2514
rect 5442 2302 5502 2416
rect 5586 2048 5646 2474
rect 5872 2474 5884 2480
rect 5924 2480 5934 2514
rect 6018 2614 6078 2630
rect 6018 2574 6028 2614
rect 6068 2574 6078 2614
rect 6018 2514 6078 2574
rect 5924 2474 5936 2480
rect 5872 2422 5878 2474
rect 5930 2422 5936 2474
rect 5872 2416 5936 2422
rect 6018 2474 6028 2514
rect 6068 2474 6078 2514
rect 6162 2614 6222 2630
rect 6162 2574 6172 2614
rect 6212 2574 6222 2614
rect 6162 2514 6222 2574
rect 6162 2480 6172 2514
rect 5874 2302 5934 2416
rect 6018 2336 6078 2474
rect 6160 2474 6172 2480
rect 6212 2480 6222 2514
rect 6450 2614 6510 2630
rect 6450 2574 6460 2614
rect 6500 2574 6510 2614
rect 6450 2514 6510 2574
rect 6212 2474 6224 2480
rect 6160 2422 6166 2474
rect 6218 2422 6224 2474
rect 6160 2416 6224 2422
rect 6450 2474 6460 2514
rect 6500 2474 6510 2514
rect 6016 2330 6080 2336
rect 6016 2278 6022 2330
rect 6074 2278 6080 2330
rect 6162 2302 6222 2416
rect 6016 2272 6080 2278
rect 5874 2048 5934 2056
rect 6162 2048 6222 2056
rect 6450 2048 6510 2474
rect 6594 2614 6654 2630
rect 6594 2574 6604 2614
rect 6644 2574 6654 2614
rect 6594 2514 6654 2574
rect 6594 2474 6604 2514
rect 6644 2474 6654 2514
rect 6594 2458 6654 2474
rect 6738 2614 6798 2630
rect 6738 2574 6748 2614
rect 6788 2574 6798 2614
rect 6738 2514 6798 2574
rect 6738 2474 6748 2514
rect 6788 2474 6798 2514
rect 6738 2336 6798 2474
rect 7026 2588 7086 2630
rect 7026 2500 7036 2588
rect 7076 2500 7086 2588
rect 6736 2330 6800 2336
rect 6736 2278 6742 2330
rect 6794 2278 6800 2330
rect 6736 2272 6800 2278
rect 6738 2048 6798 2056
rect 7026 2048 7086 2500
rect 7170 2588 7230 2630
rect 7170 2500 7180 2588
rect 7220 2500 7230 2588
rect 7170 2480 7230 2500
rect 7314 2588 7374 2630
rect 7314 2500 7324 2588
rect 7364 2500 7374 2588
rect 7168 2474 7232 2480
rect 7168 2422 7174 2474
rect 7226 2422 7232 2474
rect 7168 2416 7232 2422
rect 7170 2302 7230 2416
rect 7314 2048 7374 2500
rect 7602 2614 7662 2630
rect 7602 2574 7612 2614
rect 7652 2574 7662 2614
rect 7602 2514 7662 2574
rect 7602 2474 7612 2514
rect 7652 2474 7662 2514
rect 7746 2614 7806 2630
rect 7746 2574 7756 2614
rect 7796 2574 7806 2614
rect 7746 2514 7806 2574
rect 7746 2480 7756 2514
rect 7602 2048 7662 2474
rect 7744 2474 7756 2480
rect 7796 2480 7806 2514
rect 7890 2614 7950 2630
rect 7890 2574 7900 2614
rect 7940 2574 7950 2614
rect 7890 2514 7950 2574
rect 7796 2474 7808 2480
rect 7744 2422 7750 2474
rect 7802 2422 7808 2474
rect 7744 2416 7808 2422
rect 7890 2474 7900 2514
rect 7940 2474 7950 2514
rect 7746 2302 7806 2416
rect 7890 2048 7950 2474
rect 8178 2614 8238 2630
rect 8178 2574 8188 2614
rect 8228 2574 8238 2614
rect 8178 2514 8238 2574
rect 8178 2474 8188 2514
rect 8228 2474 8238 2514
rect 8322 2614 8382 2630
rect 8322 2574 8332 2614
rect 8372 2574 8382 2614
rect 8322 2514 8382 2574
rect 8322 2480 8332 2514
rect 8178 2048 8238 2474
rect 8320 2474 8332 2480
rect 8372 2480 8382 2514
rect 8466 2614 8526 2630
rect 8466 2574 8476 2614
rect 8516 2574 8526 2614
rect 8466 2514 8526 2574
rect 8372 2474 8384 2480
rect 8320 2422 8326 2474
rect 8378 2422 8384 2474
rect 8320 2416 8384 2422
rect 8466 2474 8476 2514
rect 8516 2474 8526 2514
rect 8754 2614 8814 2630
rect 8754 2574 8764 2614
rect 8804 2574 8814 2614
rect 8754 2514 8814 2574
rect 8754 2480 8764 2514
rect 8322 2302 8382 2416
rect 8466 2048 8526 2474
rect 8752 2474 8764 2480
rect 8804 2480 8814 2514
rect 8898 2614 8958 2630
rect 8898 2574 8908 2614
rect 8948 2574 8958 2614
rect 8898 2514 8958 2574
rect 8804 2474 8816 2480
rect 8752 2422 8758 2474
rect 8810 2422 8816 2474
rect 8752 2416 8816 2422
rect 8898 2474 8908 2514
rect 8948 2474 8958 2514
rect 9042 2614 9102 2630
rect 9042 2574 9052 2614
rect 9092 2574 9102 2614
rect 9042 2514 9102 2574
rect 9042 2480 9052 2514
rect 8754 2302 8814 2416
rect 8898 2336 8958 2474
rect 9040 2474 9052 2480
rect 9092 2480 9102 2514
rect 9330 2614 9390 2630
rect 9330 2574 9340 2614
rect 9380 2574 9390 2614
rect 9330 2514 9390 2574
rect 9092 2474 9104 2480
rect 9040 2422 9046 2474
rect 9098 2422 9104 2474
rect 9040 2416 9104 2422
rect 9330 2474 9340 2514
rect 9380 2474 9390 2514
rect 8896 2330 8960 2336
rect 8896 2278 8902 2330
rect 8954 2278 8960 2330
rect 9042 2302 9102 2416
rect 8896 2272 8960 2278
rect 8754 2048 8814 2056
rect 9042 2048 9102 2056
rect 9330 2048 9390 2474
rect 9474 2614 9534 2630
rect 9474 2574 9484 2614
rect 9524 2574 9534 2614
rect 9474 2514 9534 2574
rect 9474 2474 9484 2514
rect 9524 2474 9534 2514
rect 9474 2458 9534 2474
rect 9618 2614 9678 2630
rect 9618 2574 9628 2614
rect 9668 2574 9678 2614
rect 9618 2514 9678 2574
rect 9618 2474 9628 2514
rect 9668 2474 9678 2514
rect 9618 2336 9678 2474
rect 10194 2614 10254 2630
rect 10194 2574 10204 2614
rect 10244 2574 10254 2614
rect 10194 2514 10254 2574
rect 10194 2474 10204 2514
rect 10244 2474 10254 2514
rect 10338 2614 10398 2630
rect 10338 2574 10348 2614
rect 10388 2574 10398 2614
rect 10338 2514 10398 2574
rect 10338 2480 10348 2514
rect 9616 2330 9680 2336
rect 9616 2278 9622 2330
rect 9674 2278 9680 2330
rect 9616 2272 9680 2278
rect 9618 2048 9678 2056
rect 9906 2048 9966 2056
rect 10194 2048 10254 2474
rect 10336 2474 10348 2480
rect 10388 2480 10398 2514
rect 10482 2614 10542 2630
rect 10482 2574 10492 2614
rect 10532 2574 10542 2614
rect 10482 2514 10542 2574
rect 10388 2474 10400 2480
rect 10336 2422 10342 2474
rect 10394 2422 10400 2474
rect 10336 2416 10400 2422
rect 10482 2474 10492 2514
rect 10532 2474 10542 2514
rect 10338 2302 10398 2416
rect 10482 2048 10542 2474
rect 10770 2614 10830 2630
rect 10770 2574 10780 2614
rect 10820 2574 10830 2614
rect 10770 2514 10830 2574
rect 10770 2474 10780 2514
rect 10820 2474 10830 2514
rect 10914 2614 10974 2630
rect 10914 2574 10924 2614
rect 10964 2574 10974 2614
rect 10914 2514 10974 2574
rect 10914 2480 10924 2514
rect 10770 2048 10830 2474
rect 10912 2474 10924 2480
rect 10964 2480 10974 2514
rect 11058 2614 11118 2630
rect 11058 2574 11068 2614
rect 11108 2574 11118 2614
rect 11058 2514 11118 2574
rect 10964 2474 10976 2480
rect 10912 2422 10918 2474
rect 10970 2422 10976 2474
rect 10912 2416 10976 2422
rect 11058 2474 11068 2514
rect 11108 2474 11118 2514
rect 10914 2302 10974 2416
rect 11058 2048 11118 2474
rect 11346 2588 11406 2630
rect 11346 2500 11356 2588
rect 11396 2500 11406 2588
rect 11346 2048 11406 2500
rect 11490 2588 11550 2630
rect 11490 2500 11500 2588
rect 11540 2500 11550 2588
rect 11490 2480 11550 2500
rect 11634 2588 11694 2630
rect 11634 2500 11644 2588
rect 11684 2500 11694 2588
rect 11488 2474 11552 2480
rect 11488 2422 11494 2474
rect 11546 2422 11552 2474
rect 11488 2416 11552 2422
rect 11490 2302 11550 2416
rect 11634 2048 11694 2500
rect 11922 2614 11982 2630
rect 11922 2574 11932 2614
rect 11972 2574 11982 2614
rect 11922 2514 11982 2574
rect 11922 2474 11932 2514
rect 11972 2474 11982 2514
rect 12066 2614 12126 2630
rect 12066 2574 12076 2614
rect 12116 2574 12126 2614
rect 12066 2514 12126 2574
rect 12066 2480 12076 2514
rect 11922 2048 11982 2474
rect 12064 2474 12076 2480
rect 12116 2480 12126 2514
rect 12210 2614 12270 2630
rect 12210 2574 12220 2614
rect 12260 2574 12270 2614
rect 12210 2514 12270 2574
rect 12116 2474 12128 2480
rect 12064 2422 12070 2474
rect 12122 2422 12128 2474
rect 12064 2416 12128 2422
rect 12210 2474 12220 2514
rect 12260 2474 12270 2514
rect 12066 2302 12126 2416
rect 12210 2048 12270 2474
rect 12498 2614 12558 2630
rect 12498 2574 12508 2614
rect 12548 2574 12558 2614
rect 12498 2514 12558 2574
rect 12498 2474 12508 2514
rect 12548 2474 12558 2514
rect 12642 2614 12702 2630
rect 12642 2574 12652 2614
rect 12692 2574 12702 2614
rect 12642 2514 12702 2574
rect 12642 2480 12652 2514
rect 12498 2336 12558 2474
rect 12640 2474 12652 2480
rect 12692 2480 12702 2514
rect 12786 2614 12846 2630
rect 12786 2574 12796 2614
rect 12836 2574 12846 2614
rect 12786 2514 12846 2574
rect 12692 2474 12704 2480
rect 12640 2422 12646 2474
rect 12698 2422 12704 2474
rect 12640 2416 12704 2422
rect 12786 2474 12796 2514
rect 12836 2474 12846 2514
rect 12496 2330 12560 2336
rect 12496 2278 12502 2330
rect 12554 2278 12560 2330
rect 12642 2302 12702 2416
rect 12786 2336 12846 2474
rect 13650 2614 13710 2630
rect 13650 2574 13660 2614
rect 13700 2574 13710 2614
rect 13650 2514 13710 2574
rect 13650 2474 13660 2514
rect 13700 2474 13710 2514
rect 13794 2614 13854 2630
rect 13794 2574 13804 2614
rect 13844 2574 13854 2614
rect 13794 2514 13854 2574
rect 13794 2480 13804 2514
rect 13650 2336 13710 2474
rect 13792 2474 13804 2480
rect 13844 2480 13854 2514
rect 13938 2614 13998 2630
rect 13938 2574 13948 2614
rect 13988 2574 13998 2614
rect 13938 2514 13998 2574
rect 13844 2474 13856 2480
rect 13792 2422 13798 2474
rect 13850 2422 13856 2474
rect 13792 2416 13856 2422
rect 13938 2474 13948 2514
rect 13988 2474 13998 2514
rect 12784 2330 12848 2336
rect 12496 2272 12560 2278
rect 12784 2278 12790 2330
rect 12842 2278 12848 2330
rect 12784 2272 12848 2278
rect 13648 2330 13712 2336
rect 13648 2278 13654 2330
rect 13706 2278 13712 2330
rect 13794 2302 13854 2416
rect 13938 2336 13998 2474
rect 14226 2614 14286 2630
rect 14226 2574 14236 2614
rect 14276 2574 14286 2614
rect 14226 2514 14286 2574
rect 14226 2474 14236 2514
rect 14276 2474 14286 2514
rect 14370 2614 14430 2630
rect 14370 2574 14380 2614
rect 14420 2574 14430 2614
rect 14370 2514 14430 2574
rect 14370 2480 14380 2514
rect 13936 2330 14000 2336
rect 13648 2272 13712 2278
rect 13936 2278 13942 2330
rect 13994 2278 14000 2330
rect 13936 2272 14000 2278
rect 12498 2048 12558 2056
rect 12786 2048 12846 2056
rect 13074 2048 13134 2056
rect 13362 2048 13422 2056
rect 13650 2048 13710 2056
rect 13938 2048 13998 2056
rect 14226 2048 14286 2474
rect 14368 2474 14380 2480
rect 14420 2480 14430 2514
rect 14514 2614 14574 2630
rect 14514 2574 14524 2614
rect 14564 2574 14574 2614
rect 14514 2514 14574 2574
rect 14420 2474 14432 2480
rect 14368 2422 14374 2474
rect 14426 2422 14432 2474
rect 14368 2416 14432 2422
rect 14514 2474 14524 2514
rect 14564 2474 14574 2514
rect 14370 2302 14430 2416
rect 14514 2048 14574 2474
rect 14802 2614 14862 2630
rect 14802 2574 14812 2614
rect 14852 2574 14862 2614
rect 14802 2514 14862 2574
rect 14802 2474 14812 2514
rect 14852 2474 14862 2514
rect 14946 2614 15006 2630
rect 14946 2574 14956 2614
rect 14996 2574 15006 2614
rect 14946 2514 15006 2574
rect 14946 2480 14956 2514
rect 14802 2048 14862 2474
rect 14944 2474 14956 2480
rect 14996 2480 15006 2514
rect 15090 2614 15150 2630
rect 15090 2574 15100 2614
rect 15140 2574 15150 2614
rect 15090 2514 15150 2574
rect 14996 2474 15008 2480
rect 14944 2422 14950 2474
rect 15002 2422 15008 2474
rect 14944 2416 15008 2422
rect 15090 2474 15100 2514
rect 15140 2474 15150 2514
rect 14946 2302 15006 2416
rect 15090 2048 15150 2474
rect 15378 2588 15438 2630
rect 15378 2500 15388 2588
rect 15428 2500 15438 2588
rect 15378 2048 15438 2500
rect 15522 2588 15582 2630
rect 15522 2500 15532 2588
rect 15572 2500 15582 2588
rect 15522 2480 15582 2500
rect 15666 2588 15726 2630
rect 15666 2500 15676 2588
rect 15716 2500 15726 2588
rect 15520 2474 15584 2480
rect 15520 2422 15526 2474
rect 15578 2422 15584 2474
rect 15520 2416 15584 2422
rect 15522 2302 15582 2416
rect 15666 2048 15726 2500
rect 15954 2588 16014 2630
rect 15954 2500 15964 2588
rect 16004 2500 16014 2588
rect 15954 2048 16014 2500
rect 16098 2588 16158 2630
rect 16098 2500 16108 2588
rect 16148 2500 16158 2588
rect 16098 2480 16158 2500
rect 16242 2588 16302 2630
rect 16242 2500 16252 2588
rect 16292 2500 16302 2588
rect 16096 2474 16160 2480
rect 16096 2422 16102 2474
rect 16154 2422 16160 2474
rect 16096 2416 16160 2422
rect 16098 2302 16158 2416
rect 16242 2048 16302 2500
rect 16530 2614 16590 2630
rect 16530 2574 16540 2614
rect 16580 2574 16590 2614
rect 16530 2514 16590 2574
rect 16530 2474 16540 2514
rect 16580 2474 16590 2514
rect 16674 2614 16734 2630
rect 16674 2574 16684 2614
rect 16724 2574 16734 2614
rect 16674 2514 16734 2574
rect 16674 2480 16684 2514
rect 16530 2048 16590 2474
rect 16672 2474 16684 2480
rect 16724 2480 16734 2514
rect 16818 2614 16878 2630
rect 16818 2574 16828 2614
rect 16868 2574 16878 2614
rect 16818 2514 16878 2574
rect 16724 2474 16736 2480
rect 16672 2422 16678 2474
rect 16730 2422 16736 2474
rect 16672 2416 16736 2422
rect 16818 2474 16828 2514
rect 16868 2474 16878 2514
rect 16962 2614 17022 2630
rect 16962 2574 16972 2614
rect 17012 2574 17022 2614
rect 16962 2514 17022 2574
rect 16962 2480 16972 2514
rect 16674 2302 16734 2416
rect 16818 2048 16878 2474
rect 16960 2474 16972 2480
rect 17012 2480 17022 2514
rect 17106 2614 17166 2630
rect 17106 2574 17116 2614
rect 17156 2574 17166 2614
rect 17106 2514 17166 2574
rect 17012 2474 17024 2480
rect 16960 2422 16966 2474
rect 17018 2422 17024 2474
rect 16960 2416 17024 2422
rect 17106 2474 17116 2514
rect 17156 2474 17166 2514
rect 17250 2614 17310 2630
rect 17250 2574 17260 2614
rect 17300 2574 17310 2614
rect 17250 2514 17310 2574
rect 17250 2480 17260 2514
rect 16962 2302 17022 2416
rect 17106 2048 17166 2474
rect 17248 2474 17260 2480
rect 17300 2480 17310 2514
rect 17394 2614 17454 2630
rect 17394 2574 17404 2614
rect 17444 2574 17454 2614
rect 17394 2514 17454 2574
rect 17300 2474 17312 2480
rect 17248 2422 17254 2474
rect 17306 2422 17312 2474
rect 17248 2416 17312 2422
rect 17394 2474 17404 2514
rect 17444 2474 17454 2514
rect 17538 2614 17598 2630
rect 17538 2574 17548 2614
rect 17588 2574 17598 2614
rect 17538 2514 17598 2574
rect 17538 2480 17548 2514
rect 17250 2302 17310 2416
rect 17394 2048 17454 2474
rect 17536 2474 17548 2480
rect 17588 2480 17598 2514
rect 17682 2614 17742 2630
rect 17682 2574 17692 2614
rect 17732 2574 17742 2614
rect 17682 2514 17742 2574
rect 17588 2474 17600 2480
rect 17536 2422 17542 2474
rect 17594 2422 17600 2474
rect 17536 2416 17600 2422
rect 17682 2474 17692 2514
rect 17732 2474 17742 2514
rect 17826 2614 17886 2630
rect 17826 2574 17836 2614
rect 17876 2574 17886 2614
rect 17826 2514 17886 2574
rect 17826 2480 17836 2514
rect 17538 2302 17598 2416
rect 17682 2048 17742 2474
rect 17824 2474 17836 2480
rect 17876 2480 17886 2514
rect 17970 2614 18030 2630
rect 17970 2574 17980 2614
rect 18020 2574 18030 2614
rect 17970 2514 18030 2574
rect 17876 2474 17888 2480
rect 17824 2422 17830 2474
rect 17882 2422 17888 2474
rect 17824 2416 17888 2422
rect 17970 2474 17980 2514
rect 18020 2474 18030 2514
rect 18114 2614 18174 2630
rect 18114 2574 18124 2614
rect 18164 2574 18174 2614
rect 18114 2514 18174 2574
rect 18114 2480 18124 2514
rect 17826 2302 17886 2416
rect 17970 2048 18030 2474
rect 18112 2474 18124 2480
rect 18164 2480 18174 2514
rect 18258 2614 18318 2630
rect 18258 2574 18268 2614
rect 18308 2574 18318 2614
rect 18258 2514 18318 2574
rect 18164 2474 18176 2480
rect 18112 2422 18118 2474
rect 18170 2422 18176 2474
rect 18112 2416 18176 2422
rect 18258 2474 18268 2514
rect 18308 2474 18318 2514
rect 18402 2614 18462 2630
rect 18402 2574 18412 2614
rect 18452 2574 18462 2614
rect 18402 2514 18462 2574
rect 18402 2480 18412 2514
rect 18114 2302 18174 2416
rect 18258 2048 18318 2474
rect 18400 2474 18412 2480
rect 18452 2480 18462 2514
rect 18546 2614 18606 2630
rect 18546 2574 18556 2614
rect 18596 2574 18606 2614
rect 18546 2514 18606 2574
rect 18452 2474 18464 2480
rect 18400 2422 18406 2474
rect 18458 2422 18464 2474
rect 18400 2416 18464 2422
rect 18546 2474 18556 2514
rect 18596 2474 18606 2514
rect 18690 2614 18750 2630
rect 18690 2574 18700 2614
rect 18740 2574 18750 2614
rect 18690 2514 18750 2574
rect 18690 2480 18700 2514
rect 18402 2302 18462 2416
rect 18546 2048 18606 2474
rect 18688 2474 18700 2480
rect 18740 2480 18750 2514
rect 18834 2614 18894 2630
rect 18834 2574 18844 2614
rect 18884 2574 18894 2614
rect 18834 2514 18894 2574
rect 18740 2474 18752 2480
rect 18688 2422 18694 2474
rect 18746 2422 18752 2474
rect 18688 2416 18752 2422
rect 18834 2474 18844 2514
rect 18884 2474 18894 2514
rect 18978 2614 19038 2630
rect 18978 2574 18988 2614
rect 19028 2574 19038 2614
rect 18978 2514 19038 2574
rect 18978 2480 18988 2514
rect 18690 2302 18750 2416
rect 18834 2048 18894 2474
rect 18976 2474 18988 2480
rect 19028 2480 19038 2514
rect 19122 2614 19182 2630
rect 19122 2574 19132 2614
rect 19172 2574 19182 2614
rect 19122 2514 19182 2574
rect 19028 2474 19040 2480
rect 18976 2422 18982 2474
rect 19034 2422 19040 2474
rect 18976 2416 19040 2422
rect 19122 2474 19132 2514
rect 19172 2474 19182 2514
rect 19266 2614 19326 2630
rect 19266 2574 19276 2614
rect 19316 2574 19326 2614
rect 19266 2514 19326 2574
rect 19266 2480 19276 2514
rect 18978 2302 19038 2416
rect 19122 2048 19182 2474
rect 19264 2474 19276 2480
rect 19316 2480 19326 2514
rect 19410 2614 19470 2630
rect 19410 2574 19420 2614
rect 19460 2574 19470 2614
rect 19410 2514 19470 2574
rect 19316 2474 19328 2480
rect 19264 2422 19270 2474
rect 19322 2422 19328 2474
rect 19264 2416 19328 2422
rect 19410 2474 19420 2514
rect 19460 2474 19470 2514
rect 19554 2614 19614 2630
rect 19554 2574 19564 2614
rect 19604 2574 19614 2614
rect 19554 2514 19614 2574
rect 19554 2480 19564 2514
rect 19266 2302 19326 2416
rect 19410 2048 19470 2474
rect 19552 2474 19564 2480
rect 19604 2480 19614 2514
rect 19698 2614 19758 2630
rect 19698 2574 19708 2614
rect 19748 2574 19758 2614
rect 19698 2514 19758 2574
rect 19604 2474 19616 2480
rect 19552 2422 19558 2474
rect 19610 2422 19616 2474
rect 19552 2416 19616 2422
rect 19698 2474 19708 2514
rect 19748 2474 19758 2514
rect 19842 2614 19902 2630
rect 19842 2574 19852 2614
rect 19892 2574 19902 2614
rect 19842 2514 19902 2574
rect 19842 2480 19852 2514
rect 19554 2302 19614 2416
rect 19698 2048 19758 2474
rect 19840 2474 19852 2480
rect 19892 2480 19902 2514
rect 19986 2614 20046 2630
rect 19986 2574 19996 2614
rect 20036 2574 20046 2614
rect 19986 2514 20046 2574
rect 19892 2474 19904 2480
rect 19840 2422 19846 2474
rect 19898 2422 19904 2474
rect 19840 2416 19904 2422
rect 19986 2474 19996 2514
rect 20036 2474 20046 2514
rect 19842 2302 19902 2416
rect 19986 2048 20046 2474
rect 20274 2048 20334 2056
rect 20562 2048 20622 2056
rect 20850 2048 20910 2056
rect 112 2042 176 2048
rect 112 1990 118 2042
rect 170 1990 176 2042
rect 112 1984 176 1990
rect 400 2042 464 2048
rect 400 1990 406 2042
rect 458 1990 464 2042
rect 400 1984 464 1990
rect 688 2042 752 2048
rect 688 1990 694 2042
rect 746 1990 752 2042
rect 688 1984 752 1990
rect 976 2042 1040 2048
rect 976 1990 982 2042
rect 1034 1990 1040 2042
rect 976 1984 1040 1990
rect 1264 2042 1328 2048
rect 1264 1990 1270 2042
rect 1322 1990 1328 2042
rect 1264 1984 1328 1990
rect 1552 2042 1616 2048
rect 1552 1990 1558 2042
rect 1610 1990 1616 2042
rect 1552 1984 1616 1990
rect 1840 2042 1904 2048
rect 1840 1990 1846 2042
rect 1898 1990 1904 2042
rect 1840 1984 1904 1990
rect 2128 2042 2192 2048
rect 2128 1990 2134 2042
rect 2186 1990 2192 2042
rect 2128 1984 2192 1990
rect 2416 2042 2480 2048
rect 2416 1990 2422 2042
rect 2474 1990 2480 2042
rect 2416 1984 2480 1990
rect 2704 2042 2768 2048
rect 2704 1990 2710 2042
rect 2762 1990 2768 2042
rect 2704 1984 2768 1990
rect 2992 2042 3056 2048
rect 2992 1990 2998 2042
rect 3050 1990 3056 2042
rect 2992 1984 3056 1990
rect 3280 2042 3344 2048
rect 3280 1990 3286 2042
rect 3338 1990 3344 2042
rect 3280 1984 3344 1990
rect 3568 2042 3632 2048
rect 3568 1990 3574 2042
rect 3626 1990 3632 2042
rect 3568 1984 3632 1990
rect 3856 2042 3920 2048
rect 3856 1990 3862 2042
rect 3914 1990 3920 2042
rect 3856 1984 3920 1990
rect 4144 2042 4208 2048
rect 4144 1990 4150 2042
rect 4202 1990 4208 2042
rect 4144 1984 4208 1990
rect 4432 2042 4496 2048
rect 4432 1990 4438 2042
rect 4490 1990 4496 2042
rect 4432 1984 4496 1990
rect 4720 2042 4784 2048
rect 4720 1990 4726 2042
rect 4778 1990 4784 2042
rect 4720 1984 4784 1990
rect 5008 2042 5072 2048
rect 5008 1990 5014 2042
rect 5066 1990 5072 2042
rect 5008 1984 5072 1990
rect 5296 2042 5360 2048
rect 5296 1990 5302 2042
rect 5354 1990 5360 2042
rect 5296 1984 5360 1990
rect 5584 2042 5648 2048
rect 5584 1990 5590 2042
rect 5642 1990 5648 2042
rect 5584 1984 5648 1990
rect 5872 2042 5936 2048
rect 5872 1990 5878 2042
rect 5930 1990 5936 2042
rect 5872 1984 5936 1990
rect 6160 2042 6224 2048
rect 6160 1990 6166 2042
rect 6218 1990 6224 2042
rect 6160 1984 6224 1990
rect 6448 2042 6512 2048
rect 6448 1990 6454 2042
rect 6506 1990 6512 2042
rect 6448 1984 6512 1990
rect 6736 2042 6800 2048
rect 6736 1990 6742 2042
rect 6794 1990 6800 2042
rect 6736 1984 6800 1990
rect 7024 2042 7088 2048
rect 7024 1990 7030 2042
rect 7082 1990 7088 2042
rect 7024 1984 7088 1990
rect 7312 2042 7376 2048
rect 7312 1990 7318 2042
rect 7370 1990 7376 2042
rect 7312 1984 7376 1990
rect 7600 2042 7664 2048
rect 7600 1990 7606 2042
rect 7658 1990 7664 2042
rect 7600 1984 7664 1990
rect 7888 2042 7952 2048
rect 7888 1990 7894 2042
rect 7946 1990 7952 2042
rect 7888 1984 7952 1990
rect 8176 2042 8240 2048
rect 8176 1990 8182 2042
rect 8234 1990 8240 2042
rect 8176 1984 8240 1990
rect 8464 2042 8528 2048
rect 8464 1990 8470 2042
rect 8522 1990 8528 2042
rect 8464 1984 8528 1990
rect 8752 2042 8816 2048
rect 8752 1990 8758 2042
rect 8810 1990 8816 2042
rect 8752 1984 8816 1990
rect 9040 2042 9104 2048
rect 9040 1990 9046 2042
rect 9098 1990 9104 2042
rect 9040 1984 9104 1990
rect 9328 2042 9392 2048
rect 9328 1990 9334 2042
rect 9386 1990 9392 2042
rect 9328 1984 9392 1990
rect 9616 2042 9680 2048
rect 9616 1990 9622 2042
rect 9674 1990 9680 2042
rect 9616 1984 9680 1990
rect 9904 2042 9968 2048
rect 9904 1990 9910 2042
rect 9962 1990 9968 2042
rect 9904 1984 9968 1990
rect 10192 2042 10256 2048
rect 10192 1990 10198 2042
rect 10250 1990 10256 2042
rect 10192 1984 10256 1990
rect 10480 2042 10544 2048
rect 10480 1990 10486 2042
rect 10538 1990 10544 2042
rect 10480 1984 10544 1990
rect 10768 2042 10832 2048
rect 10768 1990 10774 2042
rect 10826 1990 10832 2042
rect 10768 1984 10832 1990
rect 11056 2042 11120 2048
rect 11056 1990 11062 2042
rect 11114 1990 11120 2042
rect 11056 1984 11120 1990
rect 11344 2042 11408 2048
rect 11344 1990 11350 2042
rect 11402 1990 11408 2042
rect 11344 1984 11408 1990
rect 11632 2042 11696 2048
rect 11632 1990 11638 2042
rect 11690 1990 11696 2042
rect 11632 1984 11696 1990
rect 11920 2042 11984 2048
rect 11920 1990 11926 2042
rect 11978 1990 11984 2042
rect 11920 1984 11984 1990
rect 12208 2042 12272 2048
rect 12208 1990 12214 2042
rect 12266 1990 12272 2042
rect 12208 1984 12272 1990
rect 12496 2042 12560 2048
rect 12496 1990 12502 2042
rect 12554 1990 12560 2042
rect 12496 1984 12560 1990
rect 12784 2042 12848 2048
rect 12784 1990 12790 2042
rect 12842 1990 12848 2042
rect 12784 1984 12848 1990
rect 13072 2042 13136 2048
rect 13072 1990 13078 2042
rect 13130 1990 13136 2042
rect 13072 1984 13136 1990
rect 13360 2042 13424 2048
rect 13360 1990 13366 2042
rect 13418 1990 13424 2042
rect 13360 1984 13424 1990
rect 13648 2042 13712 2048
rect 13648 1990 13654 2042
rect 13706 1990 13712 2042
rect 13648 1984 13712 1990
rect 13936 2042 14000 2048
rect 13936 1990 13942 2042
rect 13994 1990 14000 2042
rect 13936 1984 14000 1990
rect 14224 2042 14288 2048
rect 14224 1990 14230 2042
rect 14282 1990 14288 2042
rect 14224 1984 14288 1990
rect 14512 2042 14576 2048
rect 14512 1990 14518 2042
rect 14570 1990 14576 2042
rect 14512 1984 14576 1990
rect 14800 2042 14864 2048
rect 14800 1990 14806 2042
rect 14858 1990 14864 2042
rect 14800 1984 14864 1990
rect 15088 2042 15152 2048
rect 15088 1990 15094 2042
rect 15146 1990 15152 2042
rect 15088 1984 15152 1990
rect 15376 2042 15440 2048
rect 15376 1990 15382 2042
rect 15434 1990 15440 2042
rect 15376 1984 15440 1990
rect 15664 2042 15728 2048
rect 15664 1990 15670 2042
rect 15722 1990 15728 2042
rect 15664 1984 15728 1990
rect 15952 2042 16016 2048
rect 15952 1990 15958 2042
rect 16010 1990 16016 2042
rect 15952 1984 16016 1990
rect 16240 2042 16304 2048
rect 16240 1990 16246 2042
rect 16298 1990 16304 2042
rect 16240 1984 16304 1990
rect 16528 2042 16592 2048
rect 16528 1990 16534 2042
rect 16586 1990 16592 2042
rect 16528 1984 16592 1990
rect 16816 2042 16880 2048
rect 16816 1990 16822 2042
rect 16874 1990 16880 2042
rect 16816 1984 16880 1990
rect 17104 2042 17168 2048
rect 17104 1990 17110 2042
rect 17162 1990 17168 2042
rect 17104 1984 17168 1990
rect 17392 2042 17456 2048
rect 17392 1990 17398 2042
rect 17450 1990 17456 2042
rect 17392 1984 17456 1990
rect 17680 2042 17744 2048
rect 17680 1990 17686 2042
rect 17738 1990 17744 2042
rect 17680 1984 17744 1990
rect 17968 2042 18032 2048
rect 17968 1990 17974 2042
rect 18026 1990 18032 2042
rect 17968 1984 18032 1990
rect 18256 2042 18320 2048
rect 18256 1990 18262 2042
rect 18314 1990 18320 2042
rect 18256 1984 18320 1990
rect 18544 2042 18608 2048
rect 18544 1990 18550 2042
rect 18602 1990 18608 2042
rect 18544 1984 18608 1990
rect 18832 2042 18896 2048
rect 18832 1990 18838 2042
rect 18890 1990 18896 2042
rect 18832 1984 18896 1990
rect 19120 2042 19184 2048
rect 19120 1990 19126 2042
rect 19178 1990 19184 2042
rect 19120 1984 19184 1990
rect 19408 2042 19472 2048
rect 19408 1990 19414 2042
rect 19466 1990 19472 2042
rect 19408 1984 19472 1990
rect 19696 2042 19760 2048
rect 19696 1990 19702 2042
rect 19754 1990 19760 2042
rect 19696 1984 19760 1990
rect 19984 2042 20048 2048
rect 19984 1990 19990 2042
rect 20042 1990 20048 2042
rect 19984 1984 20048 1990
rect 20272 2042 20336 2048
rect 20272 1990 20278 2042
rect 20330 1990 20336 2042
rect 20272 1984 20336 1990
rect 20560 2042 20624 2048
rect 20560 1990 20566 2042
rect 20618 1990 20624 2042
rect 20560 1984 20624 1990
rect 20848 2042 20912 2048
rect 20848 1990 20854 2042
rect 20906 1990 20912 2042
rect 20848 1984 20912 1990
rect 114 1532 174 1984
rect 258 1616 318 1730
rect 256 1610 320 1616
rect 256 1558 262 1610
rect 314 1558 320 1610
rect 256 1552 320 1558
rect 114 1444 124 1532
rect 164 1444 174 1532
rect 114 1402 174 1444
rect 258 1532 318 1552
rect 258 1444 268 1532
rect 308 1444 318 1532
rect 258 1402 318 1444
rect 402 1532 462 1984
rect 402 1444 412 1532
rect 452 1444 462 1532
rect 402 1402 462 1444
rect 690 1558 750 1984
rect 834 1616 894 1730
rect 690 1518 700 1558
rect 740 1518 750 1558
rect 832 1610 896 1616
rect 832 1558 838 1610
rect 890 1558 896 1610
rect 832 1552 844 1558
rect 690 1458 750 1518
rect 690 1418 700 1458
rect 740 1418 750 1458
rect 690 1402 750 1418
rect 834 1518 844 1552
rect 884 1552 896 1558
rect 978 1558 1038 1984
rect 884 1518 894 1552
rect 834 1458 894 1518
rect 834 1418 844 1458
rect 884 1418 894 1458
rect 834 1402 894 1418
rect 978 1518 988 1558
rect 1028 1518 1038 1558
rect 978 1458 1038 1518
rect 978 1418 988 1458
rect 1028 1418 1038 1458
rect 978 1402 1038 1418
rect 1266 1558 1326 1984
rect 1410 1616 1470 1730
rect 1266 1518 1276 1558
rect 1316 1518 1326 1558
rect 1408 1610 1472 1616
rect 1408 1558 1414 1610
rect 1466 1558 1472 1610
rect 1408 1552 1420 1558
rect 1266 1458 1326 1518
rect 1266 1418 1276 1458
rect 1316 1418 1326 1458
rect 1266 1402 1326 1418
rect 1410 1518 1420 1552
rect 1460 1552 1472 1558
rect 1554 1558 1614 1984
rect 1842 1976 1902 1984
rect 2130 1976 2190 1984
rect 2418 1976 2478 1984
rect 2706 1976 2766 1984
rect 2994 1976 3054 1984
rect 3282 1976 3342 1984
rect 1840 1754 1904 1760
rect 1840 1702 1846 1754
rect 1898 1702 1904 1754
rect 2128 1754 2192 1760
rect 1840 1696 1904 1702
rect 1460 1518 1470 1552
rect 1410 1458 1470 1518
rect 1410 1418 1420 1458
rect 1460 1418 1470 1458
rect 1410 1402 1470 1418
rect 1554 1518 1564 1558
rect 1604 1518 1614 1558
rect 1554 1458 1614 1518
rect 1554 1418 1564 1458
rect 1604 1418 1614 1458
rect 1554 1402 1614 1418
rect 1842 1558 1902 1696
rect 1986 1616 2046 1730
rect 2128 1702 2134 1754
rect 2186 1702 2192 1754
rect 2128 1696 2192 1702
rect 2992 1754 3056 1760
rect 2992 1702 2998 1754
rect 3050 1702 3056 1754
rect 3280 1754 3344 1760
rect 2992 1696 3056 1702
rect 1842 1518 1852 1558
rect 1892 1518 1902 1558
rect 1984 1610 2048 1616
rect 1984 1558 1990 1610
rect 2042 1558 2048 1610
rect 1984 1552 1996 1558
rect 1842 1458 1902 1518
rect 1842 1418 1852 1458
rect 1892 1418 1902 1458
rect 1842 1402 1902 1418
rect 1986 1518 1996 1552
rect 2036 1552 2048 1558
rect 2130 1558 2190 1696
rect 2036 1518 2046 1552
rect 1986 1458 2046 1518
rect 1986 1418 1996 1458
rect 2036 1418 2046 1458
rect 1986 1402 2046 1418
rect 2130 1518 2140 1558
rect 2180 1518 2190 1558
rect 2130 1458 2190 1518
rect 2130 1418 2140 1458
rect 2180 1418 2190 1458
rect 2130 1402 2190 1418
rect 2994 1558 3054 1696
rect 3138 1616 3198 1730
rect 3280 1702 3286 1754
rect 3338 1702 3344 1754
rect 3280 1696 3344 1702
rect 2994 1518 3004 1558
rect 3044 1518 3054 1558
rect 3136 1610 3200 1616
rect 3136 1558 3142 1610
rect 3194 1558 3200 1610
rect 3136 1552 3148 1558
rect 2994 1458 3054 1518
rect 2994 1418 3004 1458
rect 3044 1418 3054 1458
rect 2994 1402 3054 1418
rect 3138 1518 3148 1552
rect 3188 1552 3200 1558
rect 3282 1558 3342 1696
rect 3188 1518 3198 1552
rect 3138 1458 3198 1518
rect 3138 1418 3148 1458
rect 3188 1418 3198 1458
rect 3138 1402 3198 1418
rect 3282 1518 3292 1558
rect 3332 1518 3342 1558
rect 3282 1458 3342 1518
rect 3282 1418 3292 1458
rect 3332 1418 3342 1458
rect 3282 1402 3342 1418
rect 3570 1558 3630 1984
rect 3714 1616 3774 1730
rect 3570 1518 3580 1558
rect 3620 1518 3630 1558
rect 3712 1610 3776 1616
rect 3712 1558 3718 1610
rect 3770 1558 3776 1610
rect 3712 1552 3724 1558
rect 3570 1458 3630 1518
rect 3570 1418 3580 1458
rect 3620 1418 3630 1458
rect 3570 1402 3630 1418
rect 3714 1518 3724 1552
rect 3764 1552 3776 1558
rect 3858 1558 3918 1984
rect 3764 1518 3774 1552
rect 3714 1458 3774 1518
rect 3714 1418 3724 1458
rect 3764 1418 3774 1458
rect 3714 1402 3774 1418
rect 3858 1518 3868 1558
rect 3908 1518 3918 1558
rect 3858 1458 3918 1518
rect 3858 1418 3868 1458
rect 3908 1418 3918 1458
rect 3858 1402 3918 1418
rect 4146 1558 4206 1984
rect 4290 1616 4350 1730
rect 4146 1518 4156 1558
rect 4196 1518 4206 1558
rect 4288 1610 4352 1616
rect 4288 1558 4294 1610
rect 4346 1558 4352 1610
rect 4288 1552 4300 1558
rect 4146 1458 4206 1518
rect 4146 1418 4156 1458
rect 4196 1418 4206 1458
rect 4146 1402 4206 1418
rect 4290 1518 4300 1552
rect 4340 1552 4352 1558
rect 4434 1558 4494 1984
rect 4340 1518 4350 1552
rect 4290 1458 4350 1518
rect 4290 1418 4300 1458
rect 4340 1418 4350 1458
rect 4290 1402 4350 1418
rect 4434 1518 4444 1558
rect 4484 1518 4494 1558
rect 4434 1458 4494 1518
rect 4434 1418 4444 1458
rect 4484 1418 4494 1458
rect 4434 1402 4494 1418
rect 4722 1532 4782 1984
rect 4866 1616 4926 1730
rect 4864 1610 4928 1616
rect 4864 1558 4870 1610
rect 4922 1558 4928 1610
rect 4864 1552 4928 1558
rect 4722 1444 4732 1532
rect 4772 1444 4782 1532
rect 4722 1402 4782 1444
rect 4866 1532 4926 1552
rect 4866 1444 4876 1532
rect 4916 1444 4926 1532
rect 4866 1402 4926 1444
rect 5010 1532 5070 1984
rect 5010 1444 5020 1532
rect 5060 1444 5070 1532
rect 5010 1402 5070 1444
rect 5298 1532 5358 1984
rect 5442 1616 5502 1730
rect 5440 1610 5504 1616
rect 5440 1558 5446 1610
rect 5498 1558 5504 1610
rect 5440 1552 5504 1558
rect 5298 1444 5308 1532
rect 5348 1444 5358 1532
rect 5298 1402 5358 1444
rect 5442 1532 5502 1552
rect 5442 1444 5452 1532
rect 5492 1444 5502 1532
rect 5442 1402 5502 1444
rect 5586 1532 5646 1984
rect 5586 1444 5596 1532
rect 5636 1444 5646 1532
rect 5586 1402 5646 1444
rect 5874 1558 5934 1984
rect 6018 1616 6078 1730
rect 5874 1518 5884 1558
rect 5924 1518 5934 1558
rect 6016 1610 6080 1616
rect 6016 1558 6022 1610
rect 6074 1558 6080 1610
rect 6016 1552 6028 1558
rect 5874 1458 5934 1518
rect 5874 1418 5884 1458
rect 5924 1418 5934 1458
rect 5874 1402 5934 1418
rect 6018 1518 6028 1552
rect 6068 1552 6080 1558
rect 6162 1558 6222 1984
rect 6068 1518 6078 1552
rect 6018 1458 6078 1518
rect 6018 1418 6028 1458
rect 6068 1418 6078 1458
rect 6018 1402 6078 1418
rect 6162 1518 6172 1558
rect 6212 1518 6222 1558
rect 6162 1458 6222 1518
rect 6162 1418 6172 1458
rect 6212 1418 6222 1458
rect 6162 1402 6222 1418
rect 6450 1558 6510 1984
rect 6594 1616 6654 1730
rect 6450 1518 6460 1558
rect 6500 1518 6510 1558
rect 6592 1610 6656 1616
rect 6592 1558 6598 1610
rect 6650 1558 6656 1610
rect 6592 1552 6604 1558
rect 6450 1458 6510 1518
rect 6450 1418 6460 1458
rect 6500 1418 6510 1458
rect 6450 1402 6510 1418
rect 6594 1518 6604 1552
rect 6644 1552 6656 1558
rect 6738 1558 6798 1984
rect 6644 1518 6654 1552
rect 6594 1458 6654 1518
rect 6594 1418 6604 1458
rect 6644 1418 6654 1458
rect 6594 1402 6654 1418
rect 6738 1518 6748 1558
rect 6788 1518 6798 1558
rect 6738 1458 6798 1518
rect 6738 1418 6748 1458
rect 6788 1418 6798 1458
rect 6738 1402 6798 1418
rect 7026 1558 7086 1984
rect 7170 1616 7230 1730
rect 7026 1518 7036 1558
rect 7076 1518 7086 1558
rect 7168 1610 7232 1616
rect 7168 1558 7174 1610
rect 7226 1558 7232 1610
rect 7168 1552 7180 1558
rect 7026 1458 7086 1518
rect 7026 1418 7036 1458
rect 7076 1418 7086 1458
rect 7026 1402 7086 1418
rect 7170 1518 7180 1552
rect 7220 1552 7232 1558
rect 7314 1558 7374 1984
rect 7602 1976 7662 1984
rect 7890 1976 7950 1984
rect 7744 1754 7808 1760
rect 7602 1616 7662 1730
rect 7744 1702 7750 1754
rect 7802 1702 7808 1754
rect 7744 1696 7808 1702
rect 7220 1518 7230 1552
rect 7170 1458 7230 1518
rect 7170 1418 7180 1458
rect 7220 1418 7230 1458
rect 7170 1402 7230 1418
rect 7314 1518 7324 1558
rect 7364 1518 7374 1558
rect 7600 1610 7664 1616
rect 7600 1558 7606 1610
rect 7658 1558 7664 1610
rect 7600 1552 7612 1558
rect 7314 1458 7374 1518
rect 7314 1418 7324 1458
rect 7364 1418 7374 1458
rect 7314 1402 7374 1418
rect 7602 1518 7612 1552
rect 7652 1552 7664 1558
rect 7746 1558 7806 1696
rect 7890 1616 7950 1730
rect 7652 1518 7662 1552
rect 7602 1458 7662 1518
rect 7602 1418 7612 1458
rect 7652 1418 7662 1458
rect 7602 1402 7662 1418
rect 7746 1518 7756 1558
rect 7796 1518 7806 1558
rect 7888 1610 7952 1616
rect 7888 1558 7894 1610
rect 7946 1558 7952 1610
rect 7888 1552 7900 1558
rect 7746 1458 7806 1518
rect 7746 1418 7756 1458
rect 7796 1418 7806 1458
rect 7746 1402 7806 1418
rect 7890 1518 7900 1552
rect 7940 1552 7952 1558
rect 8178 1558 8238 1984
rect 8466 1976 8526 1984
rect 8464 1754 8528 1760
rect 8464 1702 8470 1754
rect 8522 1702 8528 1754
rect 8464 1696 8528 1702
rect 7940 1518 7950 1552
rect 7890 1458 7950 1518
rect 7890 1418 7900 1458
rect 7940 1418 7950 1458
rect 7890 1402 7950 1418
rect 8178 1518 8188 1558
rect 8228 1518 8238 1558
rect 8178 1458 8238 1518
rect 8178 1418 8188 1458
rect 8228 1418 8238 1458
rect 8178 1402 8238 1418
rect 8322 1558 8382 1574
rect 8322 1518 8332 1558
rect 8372 1518 8382 1558
rect 8322 1458 8382 1518
rect 8322 1418 8332 1458
rect 8372 1418 8382 1458
rect 8322 1402 8382 1418
rect 8466 1558 8526 1696
rect 8466 1518 8476 1558
rect 8516 1518 8526 1558
rect 8466 1458 8526 1518
rect 8466 1418 8476 1458
rect 8516 1418 8526 1458
rect 8466 1402 8526 1418
rect 8754 1532 8814 1984
rect 8898 1616 8958 1730
rect 8896 1610 8960 1616
rect 8896 1558 8902 1610
rect 8954 1558 8960 1610
rect 8896 1552 8960 1558
rect 8754 1444 8764 1532
rect 8804 1444 8814 1532
rect 8754 1402 8814 1444
rect 8898 1532 8958 1552
rect 8898 1444 8908 1532
rect 8948 1444 8958 1532
rect 8898 1402 8958 1444
rect 9042 1532 9102 1984
rect 9042 1444 9052 1532
rect 9092 1444 9102 1532
rect 9042 1402 9102 1444
rect 9330 1558 9390 1984
rect 9474 1616 9534 1730
rect 9330 1518 9340 1558
rect 9380 1518 9390 1558
rect 9472 1610 9536 1616
rect 9472 1558 9478 1610
rect 9530 1558 9536 1610
rect 9472 1552 9484 1558
rect 9330 1458 9390 1518
rect 9330 1418 9340 1458
rect 9380 1418 9390 1458
rect 9330 1402 9390 1418
rect 9474 1518 9484 1552
rect 9524 1552 9536 1558
rect 9618 1558 9678 1984
rect 9524 1518 9534 1552
rect 9474 1458 9534 1518
rect 9474 1418 9484 1458
rect 9524 1418 9534 1458
rect 9474 1402 9534 1418
rect 9618 1518 9628 1558
rect 9668 1518 9678 1558
rect 9618 1458 9678 1518
rect 9618 1418 9628 1458
rect 9668 1418 9678 1458
rect 9618 1402 9678 1418
rect 9906 1558 9966 1984
rect 10050 1616 10110 1730
rect 9906 1518 9916 1558
rect 9956 1518 9966 1558
rect 10048 1610 10112 1616
rect 10048 1558 10054 1610
rect 10106 1558 10112 1610
rect 10048 1552 10060 1558
rect 9906 1458 9966 1518
rect 9906 1418 9916 1458
rect 9956 1418 9966 1458
rect 9906 1402 9966 1418
rect 10050 1518 10060 1552
rect 10100 1552 10112 1558
rect 10194 1558 10254 1984
rect 10482 1976 10542 1984
rect 10770 1976 10830 1984
rect 10624 1754 10688 1760
rect 10482 1616 10542 1730
rect 10624 1702 10630 1754
rect 10682 1702 10688 1754
rect 10624 1696 10688 1702
rect 10100 1518 10110 1552
rect 10050 1458 10110 1518
rect 10050 1418 10060 1458
rect 10100 1418 10110 1458
rect 10050 1402 10110 1418
rect 10194 1518 10204 1558
rect 10244 1518 10254 1558
rect 10480 1610 10544 1616
rect 10480 1558 10486 1610
rect 10538 1558 10544 1610
rect 10480 1552 10492 1558
rect 10194 1458 10254 1518
rect 10194 1418 10204 1458
rect 10244 1418 10254 1458
rect 10194 1402 10254 1418
rect 10482 1518 10492 1552
rect 10532 1552 10544 1558
rect 10626 1558 10686 1696
rect 10770 1616 10830 1730
rect 10532 1518 10542 1552
rect 10482 1458 10542 1518
rect 10482 1418 10492 1458
rect 10532 1418 10542 1458
rect 10482 1402 10542 1418
rect 10626 1518 10636 1558
rect 10676 1518 10686 1558
rect 10768 1610 10832 1616
rect 10768 1558 10774 1610
rect 10826 1558 10832 1610
rect 10768 1552 10780 1558
rect 10626 1458 10686 1518
rect 10626 1418 10636 1458
rect 10676 1418 10686 1458
rect 10626 1402 10686 1418
rect 10770 1518 10780 1552
rect 10820 1552 10832 1558
rect 11058 1558 11118 1984
rect 11346 1976 11406 1984
rect 11634 1976 11694 1984
rect 11344 1754 11408 1760
rect 11344 1702 11350 1754
rect 11402 1702 11408 1754
rect 11344 1696 11408 1702
rect 10820 1518 10830 1552
rect 10770 1458 10830 1518
rect 10770 1418 10780 1458
rect 10820 1418 10830 1458
rect 10770 1402 10830 1418
rect 11058 1518 11068 1558
rect 11108 1518 11118 1558
rect 11058 1458 11118 1518
rect 11058 1418 11068 1458
rect 11108 1418 11118 1458
rect 11058 1402 11118 1418
rect 11202 1558 11262 1574
rect 11202 1518 11212 1558
rect 11252 1518 11262 1558
rect 11202 1458 11262 1518
rect 11202 1418 11212 1458
rect 11252 1418 11262 1458
rect 11202 1402 11262 1418
rect 11346 1558 11406 1696
rect 11346 1518 11356 1558
rect 11396 1518 11406 1558
rect 11346 1458 11406 1518
rect 11346 1418 11356 1458
rect 11396 1418 11406 1458
rect 11346 1402 11406 1418
rect 11922 1558 11982 1984
rect 12066 1616 12126 1730
rect 11922 1518 11932 1558
rect 11972 1518 11982 1558
rect 12064 1610 12128 1616
rect 12064 1558 12070 1610
rect 12122 1558 12128 1610
rect 12064 1552 12076 1558
rect 11922 1458 11982 1518
rect 11922 1418 11932 1458
rect 11972 1418 11982 1458
rect 11922 1402 11982 1418
rect 12066 1518 12076 1552
rect 12116 1552 12128 1558
rect 12210 1558 12270 1984
rect 12116 1518 12126 1552
rect 12066 1458 12126 1518
rect 12066 1418 12076 1458
rect 12116 1418 12126 1458
rect 12066 1402 12126 1418
rect 12210 1518 12220 1558
rect 12260 1518 12270 1558
rect 12210 1458 12270 1518
rect 12210 1418 12220 1458
rect 12260 1418 12270 1458
rect 12210 1402 12270 1418
rect 12498 1558 12558 1984
rect 12642 1616 12702 1730
rect 12498 1518 12508 1558
rect 12548 1518 12558 1558
rect 12640 1610 12704 1616
rect 12640 1558 12646 1610
rect 12698 1558 12704 1610
rect 12640 1552 12652 1558
rect 12498 1458 12558 1518
rect 12498 1418 12508 1458
rect 12548 1418 12558 1458
rect 12498 1402 12558 1418
rect 12642 1518 12652 1552
rect 12692 1552 12704 1558
rect 12786 1558 12846 1984
rect 12692 1518 12702 1552
rect 12642 1458 12702 1518
rect 12642 1418 12652 1458
rect 12692 1418 12702 1458
rect 12642 1402 12702 1418
rect 12786 1518 12796 1558
rect 12836 1518 12846 1558
rect 12786 1458 12846 1518
rect 12786 1418 12796 1458
rect 12836 1418 12846 1458
rect 12786 1402 12846 1418
rect 13074 1558 13134 1984
rect 13218 1616 13278 1730
rect 13074 1518 13084 1558
rect 13124 1518 13134 1558
rect 13216 1610 13280 1616
rect 13216 1558 13222 1610
rect 13274 1558 13280 1610
rect 13216 1552 13228 1558
rect 13074 1458 13134 1518
rect 13074 1418 13084 1458
rect 13124 1418 13134 1458
rect 13074 1402 13134 1418
rect 13218 1518 13228 1552
rect 13268 1552 13280 1558
rect 13362 1558 13422 1984
rect 13268 1518 13278 1552
rect 13218 1458 13278 1518
rect 13218 1418 13228 1458
rect 13268 1418 13278 1458
rect 13218 1402 13278 1418
rect 13362 1518 13372 1558
rect 13412 1518 13422 1558
rect 13362 1458 13422 1518
rect 13362 1418 13372 1458
rect 13412 1418 13422 1458
rect 13362 1402 13422 1418
rect 13650 1558 13710 1984
rect 13794 1616 13854 1730
rect 13650 1518 13660 1558
rect 13700 1518 13710 1558
rect 13792 1610 13856 1616
rect 13792 1558 13798 1610
rect 13850 1558 13856 1610
rect 13792 1552 13804 1558
rect 13650 1458 13710 1518
rect 13650 1418 13660 1458
rect 13700 1418 13710 1458
rect 13650 1402 13710 1418
rect 13794 1518 13804 1552
rect 13844 1552 13856 1558
rect 13938 1558 13998 1984
rect 13844 1518 13854 1552
rect 13794 1458 13854 1518
rect 13794 1418 13804 1458
rect 13844 1418 13854 1458
rect 13794 1402 13854 1418
rect 13938 1518 13948 1558
rect 13988 1518 13998 1558
rect 13938 1458 13998 1518
rect 13938 1418 13948 1458
rect 13988 1418 13998 1458
rect 13938 1402 13998 1418
rect 14226 1532 14286 1984
rect 14370 1616 14430 1730
rect 14368 1610 14432 1616
rect 14368 1558 14374 1610
rect 14426 1558 14432 1610
rect 14368 1552 14432 1558
rect 14226 1444 14236 1532
rect 14276 1444 14286 1532
rect 14226 1402 14286 1444
rect 14370 1532 14430 1552
rect 14370 1444 14380 1532
rect 14420 1444 14430 1532
rect 14370 1402 14430 1444
rect 14514 1532 14574 1984
rect 14514 1444 14524 1532
rect 14564 1444 14574 1532
rect 14514 1402 14574 1444
rect 14802 1558 14862 1984
rect 14946 1616 15006 1730
rect 14802 1518 14812 1558
rect 14852 1518 14862 1558
rect 14944 1610 15008 1616
rect 14944 1558 14950 1610
rect 15002 1558 15008 1610
rect 14944 1552 14956 1558
rect 14802 1458 14862 1518
rect 14802 1418 14812 1458
rect 14852 1418 14862 1458
rect 14802 1402 14862 1418
rect 14946 1518 14956 1552
rect 14996 1552 15008 1558
rect 15090 1558 15150 1984
rect 14996 1518 15006 1552
rect 14946 1458 15006 1518
rect 14946 1418 14956 1458
rect 14996 1418 15006 1458
rect 14946 1402 15006 1418
rect 15090 1518 15100 1558
rect 15140 1518 15150 1558
rect 15090 1458 15150 1518
rect 15090 1418 15100 1458
rect 15140 1418 15150 1458
rect 15090 1402 15150 1418
rect 15378 1558 15438 1984
rect 15522 1616 15582 1730
rect 15378 1518 15388 1558
rect 15428 1518 15438 1558
rect 15520 1610 15584 1616
rect 15520 1558 15526 1610
rect 15578 1558 15584 1610
rect 15520 1552 15532 1558
rect 15378 1458 15438 1518
rect 15378 1418 15388 1458
rect 15428 1418 15438 1458
rect 15378 1402 15438 1418
rect 15522 1518 15532 1552
rect 15572 1552 15584 1558
rect 15666 1558 15726 1984
rect 15572 1518 15582 1552
rect 15522 1458 15582 1518
rect 15522 1418 15532 1458
rect 15572 1418 15582 1458
rect 15522 1402 15582 1418
rect 15666 1518 15676 1558
rect 15716 1518 15726 1558
rect 15666 1458 15726 1518
rect 15666 1418 15676 1458
rect 15716 1418 15726 1458
rect 15666 1402 15726 1418
rect 15954 1558 16014 1984
rect 16098 1616 16158 1730
rect 15954 1518 15964 1558
rect 16004 1518 16014 1558
rect 16096 1610 16160 1616
rect 16096 1558 16102 1610
rect 16154 1558 16160 1610
rect 16096 1552 16108 1558
rect 15954 1458 16014 1518
rect 15954 1418 15964 1458
rect 16004 1418 16014 1458
rect 15954 1402 16014 1418
rect 16098 1518 16108 1552
rect 16148 1552 16160 1558
rect 16242 1558 16302 1984
rect 16386 1616 16446 1730
rect 16148 1518 16158 1552
rect 16098 1458 16158 1518
rect 16098 1418 16108 1458
rect 16148 1418 16158 1458
rect 16098 1402 16158 1418
rect 16242 1518 16252 1558
rect 16292 1518 16302 1558
rect 16384 1610 16448 1616
rect 16384 1558 16390 1610
rect 16442 1558 16448 1610
rect 16384 1552 16396 1558
rect 16242 1458 16302 1518
rect 16242 1418 16252 1458
rect 16292 1418 16302 1458
rect 16242 1402 16302 1418
rect 16386 1518 16396 1552
rect 16436 1552 16448 1558
rect 16530 1558 16590 1984
rect 16436 1518 16446 1552
rect 16386 1458 16446 1518
rect 16386 1418 16396 1458
rect 16436 1418 16446 1458
rect 16386 1402 16446 1418
rect 16530 1518 16540 1558
rect 16580 1518 16590 1558
rect 16530 1458 16590 1518
rect 16530 1418 16540 1458
rect 16580 1418 16590 1458
rect 16530 1402 16590 1418
rect 16818 1532 16878 1984
rect 16962 1616 17022 1730
rect 16960 1610 17024 1616
rect 16960 1558 16966 1610
rect 17018 1558 17024 1610
rect 16960 1552 17024 1558
rect 16818 1444 16828 1532
rect 16868 1444 16878 1532
rect 16818 1402 16878 1444
rect 16962 1532 17022 1552
rect 16962 1444 16972 1532
rect 17012 1444 17022 1532
rect 16962 1402 17022 1444
rect 17106 1532 17166 1984
rect 17106 1444 17116 1532
rect 17156 1444 17166 1532
rect 17106 1402 17166 1444
rect 17394 1558 17454 1984
rect 17538 1616 17598 1730
rect 17394 1518 17404 1558
rect 17444 1518 17454 1558
rect 17536 1610 17600 1616
rect 17536 1558 17542 1610
rect 17594 1558 17600 1610
rect 17536 1552 17548 1558
rect 17394 1458 17454 1518
rect 17394 1418 17404 1458
rect 17444 1418 17454 1458
rect 17394 1402 17454 1418
rect 17538 1518 17548 1552
rect 17588 1552 17600 1558
rect 17682 1558 17742 1984
rect 17826 1616 17886 1730
rect 17588 1518 17598 1552
rect 17538 1458 17598 1518
rect 17538 1418 17548 1458
rect 17588 1418 17598 1458
rect 17538 1402 17598 1418
rect 17682 1518 17692 1558
rect 17732 1518 17742 1558
rect 17824 1610 17888 1616
rect 17824 1558 17830 1610
rect 17882 1558 17888 1610
rect 17824 1552 17836 1558
rect 17682 1458 17742 1518
rect 17682 1418 17692 1458
rect 17732 1418 17742 1458
rect 17682 1402 17742 1418
rect 17826 1518 17836 1552
rect 17876 1552 17888 1558
rect 17970 1558 18030 1984
rect 18114 1616 18174 1730
rect 17876 1518 17886 1552
rect 17826 1458 17886 1518
rect 17826 1418 17836 1458
rect 17876 1418 17886 1458
rect 17826 1402 17886 1418
rect 17970 1518 17980 1558
rect 18020 1518 18030 1558
rect 18112 1610 18176 1616
rect 18112 1558 18118 1610
rect 18170 1558 18176 1610
rect 18112 1552 18124 1558
rect 17970 1458 18030 1518
rect 17970 1418 17980 1458
rect 18020 1418 18030 1458
rect 17970 1402 18030 1418
rect 18114 1518 18124 1552
rect 18164 1552 18176 1558
rect 18258 1558 18318 1984
rect 18402 1616 18462 1730
rect 18164 1518 18174 1552
rect 18114 1458 18174 1518
rect 18114 1418 18124 1458
rect 18164 1418 18174 1458
rect 18114 1402 18174 1418
rect 18258 1518 18268 1558
rect 18308 1518 18318 1558
rect 18400 1610 18464 1616
rect 18400 1558 18406 1610
rect 18458 1558 18464 1610
rect 18400 1552 18412 1558
rect 18258 1458 18318 1518
rect 18258 1418 18268 1458
rect 18308 1418 18318 1458
rect 18258 1402 18318 1418
rect 18402 1518 18412 1552
rect 18452 1552 18464 1558
rect 18546 1558 18606 1984
rect 18690 1616 18750 1730
rect 18452 1518 18462 1552
rect 18402 1458 18462 1518
rect 18402 1418 18412 1458
rect 18452 1418 18462 1458
rect 18402 1402 18462 1418
rect 18546 1518 18556 1558
rect 18596 1518 18606 1558
rect 18688 1610 18752 1616
rect 18688 1558 18694 1610
rect 18746 1558 18752 1610
rect 18688 1552 18700 1558
rect 18546 1458 18606 1518
rect 18546 1418 18556 1458
rect 18596 1418 18606 1458
rect 18546 1402 18606 1418
rect 18690 1518 18700 1552
rect 18740 1552 18752 1558
rect 18834 1558 18894 1984
rect 18978 1616 19038 1730
rect 18740 1518 18750 1552
rect 18690 1458 18750 1518
rect 18690 1418 18700 1458
rect 18740 1418 18750 1458
rect 18690 1402 18750 1418
rect 18834 1518 18844 1558
rect 18884 1518 18894 1558
rect 18976 1610 19040 1616
rect 18976 1558 18982 1610
rect 19034 1558 19040 1610
rect 18976 1552 18988 1558
rect 18834 1458 18894 1518
rect 18834 1418 18844 1458
rect 18884 1418 18894 1458
rect 18834 1402 18894 1418
rect 18978 1518 18988 1552
rect 19028 1552 19040 1558
rect 19122 1558 19182 1984
rect 19266 1616 19326 1730
rect 19028 1518 19038 1552
rect 18978 1458 19038 1518
rect 18978 1418 18988 1458
rect 19028 1418 19038 1458
rect 18978 1402 19038 1418
rect 19122 1518 19132 1558
rect 19172 1518 19182 1558
rect 19264 1610 19328 1616
rect 19264 1558 19270 1610
rect 19322 1558 19328 1610
rect 19264 1552 19276 1558
rect 19122 1458 19182 1518
rect 19122 1418 19132 1458
rect 19172 1418 19182 1458
rect 19122 1402 19182 1418
rect 19266 1518 19276 1552
rect 19316 1552 19328 1558
rect 19410 1558 19470 1984
rect 19554 1616 19614 1730
rect 19316 1518 19326 1552
rect 19266 1458 19326 1518
rect 19266 1418 19276 1458
rect 19316 1418 19326 1458
rect 19266 1402 19326 1418
rect 19410 1518 19420 1558
rect 19460 1518 19470 1558
rect 19552 1610 19616 1616
rect 19552 1558 19558 1610
rect 19610 1558 19616 1610
rect 19552 1552 19564 1558
rect 19410 1458 19470 1518
rect 19410 1418 19420 1458
rect 19460 1418 19470 1458
rect 19410 1402 19470 1418
rect 19554 1518 19564 1552
rect 19604 1552 19616 1558
rect 19698 1558 19758 1984
rect 19842 1616 19902 1730
rect 19604 1518 19614 1552
rect 19554 1458 19614 1518
rect 19554 1418 19564 1458
rect 19604 1418 19614 1458
rect 19554 1402 19614 1418
rect 19698 1518 19708 1558
rect 19748 1518 19758 1558
rect 19840 1610 19904 1616
rect 19840 1558 19846 1610
rect 19898 1558 19904 1610
rect 19840 1552 19852 1558
rect 19698 1458 19758 1518
rect 19698 1418 19708 1458
rect 19748 1418 19758 1458
rect 19698 1402 19758 1418
rect 19842 1518 19852 1552
rect 19892 1552 19904 1558
rect 19986 1558 20046 1984
rect 20130 1616 20190 1730
rect 19892 1518 19902 1552
rect 19842 1458 19902 1518
rect 19842 1418 19852 1458
rect 19892 1418 19902 1458
rect 19842 1402 19902 1418
rect 19986 1518 19996 1558
rect 20036 1518 20046 1558
rect 20128 1610 20192 1616
rect 20128 1558 20134 1610
rect 20186 1558 20192 1610
rect 20128 1552 20140 1558
rect 19986 1458 20046 1518
rect 19986 1418 19996 1458
rect 20036 1418 20046 1458
rect 19986 1402 20046 1418
rect 20130 1518 20140 1552
rect 20180 1552 20192 1558
rect 20274 1558 20334 1984
rect 20418 1616 20478 1730
rect 20180 1518 20190 1552
rect 20130 1458 20190 1518
rect 20130 1418 20140 1458
rect 20180 1418 20190 1458
rect 20130 1402 20190 1418
rect 20274 1518 20284 1558
rect 20324 1518 20334 1558
rect 20416 1610 20480 1616
rect 20416 1558 20422 1610
rect 20474 1558 20480 1610
rect 20416 1552 20428 1558
rect 20274 1458 20334 1518
rect 20274 1418 20284 1458
rect 20324 1418 20334 1458
rect 20274 1402 20334 1418
rect 20418 1518 20428 1552
rect 20468 1552 20480 1558
rect 20562 1558 20622 1984
rect 20706 1616 20766 1730
rect 20468 1518 20478 1552
rect 20418 1458 20478 1518
rect 20418 1418 20428 1458
rect 20468 1418 20478 1458
rect 20418 1402 20478 1418
rect 20562 1518 20572 1558
rect 20612 1518 20622 1558
rect 20704 1610 20768 1616
rect 20704 1558 20710 1610
rect 20762 1558 20768 1610
rect 20704 1552 20716 1558
rect 20562 1458 20622 1518
rect 20562 1418 20572 1458
rect 20612 1418 20622 1458
rect 20562 1402 20622 1418
rect 20706 1518 20716 1552
rect 20756 1552 20768 1558
rect 20850 1558 20910 1984
rect 20756 1518 20766 1552
rect 20706 1458 20766 1518
rect 20706 1418 20716 1458
rect 20756 1418 20766 1458
rect 20706 1402 20766 1418
rect 20850 1518 20860 1558
rect 20900 1518 20910 1558
rect 20850 1458 20910 1518
rect 20850 1418 20860 1458
rect 20900 1418 20910 1458
rect 20850 1402 20910 1418
rect 776 1322 950 1332
rect 776 1313 838 1322
rect 776 1279 796 1313
rect 830 1279 838 1313
rect 776 1270 838 1279
rect 890 1313 950 1322
rect 890 1279 904 1313
rect 938 1279 950 1313
rect 890 1270 950 1279
rect 776 1260 950 1270
rect 1352 1322 1526 1332
rect 1352 1313 1414 1322
rect 1352 1279 1372 1313
rect 1406 1279 1414 1313
rect 1352 1270 1414 1279
rect 1466 1313 1526 1322
rect 1466 1279 1480 1313
rect 1514 1279 1526 1313
rect 1466 1270 1526 1279
rect 1352 1260 1526 1270
rect 1928 1322 2102 1332
rect 1928 1313 1990 1322
rect 1928 1279 1948 1313
rect 1982 1279 1990 1313
rect 1928 1270 1990 1279
rect 2042 1313 2102 1322
rect 2042 1279 2056 1313
rect 2090 1279 2102 1313
rect 2042 1270 2102 1279
rect 1928 1260 2102 1270
rect 3080 1322 3254 1332
rect 3080 1313 3142 1322
rect 3080 1279 3100 1313
rect 3134 1279 3142 1313
rect 3080 1270 3142 1279
rect 3194 1313 3254 1322
rect 3194 1279 3208 1313
rect 3242 1279 3254 1313
rect 3194 1270 3254 1279
rect 3080 1260 3254 1270
rect 3656 1322 3830 1332
rect 3656 1313 3718 1322
rect 3656 1279 3676 1313
rect 3710 1279 3718 1313
rect 3656 1270 3718 1279
rect 3770 1313 3830 1322
rect 3770 1279 3784 1313
rect 3818 1279 3830 1313
rect 3770 1270 3830 1279
rect 3656 1260 3830 1270
rect 4232 1322 4406 1332
rect 4232 1313 4294 1322
rect 4232 1279 4252 1313
rect 4286 1279 4294 1313
rect 4232 1270 4294 1279
rect 4346 1313 4406 1322
rect 4346 1279 4360 1313
rect 4394 1279 4406 1313
rect 4346 1270 4406 1279
rect 4232 1260 4406 1270
rect 5960 1322 6134 1332
rect 5960 1313 6022 1322
rect 5960 1279 5980 1313
rect 6014 1279 6022 1313
rect 5960 1270 6022 1279
rect 6074 1313 6134 1322
rect 6074 1279 6088 1313
rect 6122 1279 6134 1313
rect 6074 1270 6134 1279
rect 5960 1260 6134 1270
rect 6536 1322 6710 1332
rect 6536 1313 6598 1322
rect 6536 1279 6556 1313
rect 6590 1279 6598 1313
rect 6536 1270 6598 1279
rect 6650 1313 6710 1322
rect 6650 1279 6664 1313
rect 6698 1279 6710 1313
rect 6650 1270 6710 1279
rect 6536 1260 6710 1270
rect 7112 1322 7286 1332
rect 7112 1313 7174 1322
rect 7112 1279 7132 1313
rect 7166 1279 7174 1313
rect 7112 1270 7174 1279
rect 7226 1313 7286 1322
rect 7226 1279 7240 1313
rect 7274 1279 7286 1313
rect 7226 1270 7286 1279
rect 7112 1260 7286 1270
rect 7688 1322 7862 1332
rect 7688 1313 7750 1322
rect 7688 1279 7708 1313
rect 7742 1279 7750 1313
rect 7688 1270 7750 1279
rect 7802 1313 7862 1322
rect 7802 1279 7816 1313
rect 7850 1279 7862 1313
rect 7802 1270 7862 1279
rect 7688 1260 7862 1270
rect 8174 1314 8264 1332
rect 8174 1278 8196 1314
rect 8232 1278 8264 1314
rect 8174 1260 8264 1278
rect 8438 1322 8528 1332
rect 8438 1270 8470 1322
rect 8522 1270 8528 1322
rect 8438 1260 8528 1270
rect 9416 1322 9590 1332
rect 9416 1313 9478 1322
rect 9416 1279 9436 1313
rect 9470 1279 9478 1313
rect 9416 1270 9478 1279
rect 9530 1313 9590 1322
rect 9530 1279 9544 1313
rect 9578 1279 9590 1313
rect 9530 1270 9590 1279
rect 9416 1260 9590 1270
rect 9992 1322 10166 1332
rect 9992 1313 10054 1322
rect 9992 1279 10012 1313
rect 10046 1279 10054 1313
rect 9992 1270 10054 1279
rect 10106 1313 10166 1322
rect 10106 1279 10120 1313
rect 10154 1279 10166 1313
rect 10106 1270 10166 1279
rect 9992 1260 10166 1270
rect 10568 1322 10742 1332
rect 10568 1313 10630 1322
rect 10568 1279 10588 1313
rect 10622 1279 10630 1313
rect 10568 1270 10630 1279
rect 10682 1313 10742 1322
rect 10682 1279 10696 1313
rect 10730 1279 10742 1313
rect 10682 1270 10742 1279
rect 10568 1260 10742 1270
rect 11054 1314 11144 1332
rect 11054 1278 11076 1314
rect 11112 1278 11144 1314
rect 11054 1260 11144 1278
rect 11318 1322 11408 1332
rect 11318 1270 11350 1322
rect 11402 1270 11408 1322
rect 11318 1260 11408 1270
rect 12008 1322 12182 1332
rect 12008 1313 12070 1322
rect 12008 1279 12028 1313
rect 12062 1279 12070 1313
rect 12008 1270 12070 1279
rect 12122 1313 12182 1322
rect 12122 1279 12136 1313
rect 12170 1279 12182 1313
rect 12122 1270 12182 1279
rect 12008 1260 12182 1270
rect 12584 1322 12758 1332
rect 12584 1313 12646 1322
rect 12584 1279 12604 1313
rect 12638 1279 12646 1313
rect 12584 1270 12646 1279
rect 12698 1313 12758 1322
rect 12698 1279 12712 1313
rect 12746 1279 12758 1313
rect 12698 1270 12758 1279
rect 12584 1260 12758 1270
rect 13160 1322 13334 1332
rect 13160 1313 13222 1322
rect 13160 1279 13180 1313
rect 13214 1279 13222 1313
rect 13160 1270 13222 1279
rect 13274 1313 13334 1322
rect 13274 1279 13288 1313
rect 13322 1279 13334 1313
rect 13274 1270 13334 1279
rect 13160 1260 13334 1270
rect 13736 1322 13910 1332
rect 13736 1313 13798 1322
rect 13736 1279 13756 1313
rect 13790 1279 13798 1313
rect 13736 1270 13798 1279
rect 13850 1313 13910 1322
rect 13850 1279 13864 1313
rect 13898 1279 13910 1313
rect 13850 1270 13910 1279
rect 13736 1260 13910 1270
rect 14888 1322 15062 1332
rect 14888 1313 14950 1322
rect 14888 1279 14908 1313
rect 14942 1279 14950 1313
rect 14888 1270 14950 1279
rect 15002 1313 15062 1322
rect 15002 1279 15016 1313
rect 15050 1279 15062 1313
rect 15002 1270 15062 1279
rect 14888 1260 15062 1270
rect 15466 1322 15640 1332
rect 15466 1313 15526 1322
rect 15466 1279 15478 1313
rect 15512 1279 15526 1313
rect 15466 1270 15526 1279
rect 15578 1313 15640 1322
rect 15578 1279 15586 1313
rect 15620 1279 15640 1313
rect 15578 1270 15640 1279
rect 15466 1260 15640 1270
rect 16040 1322 16214 1332
rect 16040 1313 16102 1322
rect 16040 1279 16060 1313
rect 16094 1279 16102 1313
rect 16040 1270 16102 1279
rect 16154 1313 16214 1322
rect 16154 1279 16168 1313
rect 16202 1279 16214 1313
rect 16154 1270 16214 1279
rect 16040 1260 16214 1270
rect 16328 1322 16502 1332
rect 16328 1313 16390 1322
rect 16328 1279 16348 1313
rect 16382 1279 16390 1313
rect 16328 1270 16390 1279
rect 16442 1313 16502 1322
rect 16442 1279 16456 1313
rect 16490 1279 16502 1313
rect 16442 1270 16502 1279
rect 16328 1260 16502 1270
rect 17480 1322 17654 1332
rect 17480 1313 17542 1322
rect 17480 1279 17500 1313
rect 17534 1279 17542 1313
rect 17480 1270 17542 1279
rect 17594 1313 17654 1322
rect 17594 1279 17608 1313
rect 17642 1279 17654 1313
rect 17594 1270 17654 1279
rect 17480 1260 17654 1270
rect 17768 1322 17942 1332
rect 17768 1313 17830 1322
rect 17768 1279 17788 1313
rect 17822 1279 17830 1313
rect 17768 1270 17830 1279
rect 17882 1313 17942 1322
rect 17882 1279 17896 1313
rect 17930 1279 17942 1313
rect 17882 1270 17942 1279
rect 17768 1260 17942 1270
rect 18056 1322 18230 1332
rect 18056 1313 18118 1322
rect 18056 1279 18076 1313
rect 18110 1279 18118 1313
rect 18056 1270 18118 1279
rect 18170 1313 18230 1322
rect 18170 1279 18184 1313
rect 18218 1279 18230 1313
rect 18170 1270 18230 1279
rect 18056 1260 18230 1270
rect 18344 1322 18518 1332
rect 18344 1313 18406 1322
rect 18344 1279 18364 1313
rect 18398 1279 18406 1313
rect 18344 1270 18406 1279
rect 18458 1313 18518 1322
rect 18458 1279 18472 1313
rect 18506 1279 18518 1313
rect 18458 1270 18518 1279
rect 18344 1260 18518 1270
rect 18632 1322 18806 1332
rect 18632 1313 18694 1322
rect 18632 1279 18652 1313
rect 18686 1279 18694 1313
rect 18632 1270 18694 1279
rect 18746 1313 18806 1322
rect 18746 1279 18760 1313
rect 18794 1279 18806 1313
rect 18746 1270 18806 1279
rect 18632 1260 18806 1270
rect 18920 1322 19094 1332
rect 18920 1313 18982 1322
rect 18920 1279 18940 1313
rect 18974 1279 18982 1313
rect 18920 1270 18982 1279
rect 19034 1313 19094 1322
rect 19034 1279 19048 1313
rect 19082 1279 19094 1313
rect 19034 1270 19094 1279
rect 18920 1260 19094 1270
rect 19208 1322 19382 1332
rect 19208 1313 19270 1322
rect 19208 1279 19228 1313
rect 19262 1279 19270 1313
rect 19208 1270 19270 1279
rect 19322 1313 19382 1322
rect 19322 1279 19336 1313
rect 19370 1279 19382 1313
rect 19322 1270 19382 1279
rect 19208 1260 19382 1270
rect 19496 1322 19670 1332
rect 19496 1313 19558 1322
rect 19496 1279 19516 1313
rect 19550 1279 19558 1313
rect 19496 1270 19558 1279
rect 19610 1313 19670 1322
rect 19610 1279 19624 1313
rect 19658 1279 19670 1313
rect 19610 1270 19670 1279
rect 19496 1260 19670 1270
rect 19784 1322 19958 1332
rect 19784 1313 19846 1322
rect 19784 1279 19804 1313
rect 19838 1279 19846 1313
rect 19784 1270 19846 1279
rect 19898 1313 19958 1322
rect 19898 1279 19912 1313
rect 19946 1279 19958 1313
rect 19898 1270 19958 1279
rect 19784 1260 19958 1270
rect 20072 1322 20246 1332
rect 20072 1313 20134 1322
rect 20072 1279 20092 1313
rect 20126 1279 20134 1313
rect 20072 1270 20134 1279
rect 20186 1313 20246 1322
rect 20186 1279 20200 1313
rect 20234 1279 20246 1313
rect 20186 1270 20246 1279
rect 20072 1260 20246 1270
rect 20360 1322 20534 1332
rect 20360 1313 20422 1322
rect 20360 1279 20380 1313
rect 20414 1279 20422 1313
rect 20360 1270 20422 1279
rect 20474 1313 20534 1322
rect 20474 1279 20488 1313
rect 20522 1279 20534 1313
rect 20474 1270 20534 1279
rect 20360 1260 20534 1270
rect 20648 1322 20822 1332
rect 20648 1313 20710 1322
rect 20648 1279 20668 1313
rect 20702 1279 20710 1313
rect 20648 1270 20710 1279
rect 20762 1313 20822 1322
rect 20762 1279 20776 1313
rect 20810 1279 20822 1313
rect 20762 1270 20822 1279
rect 20648 1260 20822 1270
rect 8178 1040 8238 1260
rect 11058 1040 11118 1260
rect 8176 1034 8240 1040
rect 8176 982 8182 1034
rect 8234 982 8240 1034
rect 8176 976 8240 982
rect 11056 1034 11120 1040
rect 11056 982 11062 1034
rect 11114 982 11120 1034
rect 11056 976 11120 982
rect 8178 756 8238 976
rect 11058 756 11118 976
rect 776 746 950 756
rect 776 737 838 746
rect 776 703 796 737
rect 830 703 838 737
rect 776 694 838 703
rect 890 737 950 746
rect 890 703 904 737
rect 938 703 950 737
rect 890 694 950 703
rect 776 684 950 694
rect 1352 746 1526 756
rect 1352 737 1414 746
rect 1352 703 1372 737
rect 1406 703 1414 737
rect 1352 694 1414 703
rect 1466 737 1526 746
rect 1466 703 1480 737
rect 1514 703 1526 737
rect 1466 694 1526 703
rect 1352 684 1526 694
rect 1928 746 2102 756
rect 1928 737 1990 746
rect 1928 703 1948 737
rect 1982 703 1990 737
rect 1928 694 1990 703
rect 2042 737 2102 746
rect 2042 703 2056 737
rect 2090 703 2102 737
rect 2042 694 2102 703
rect 1928 684 2102 694
rect 3080 746 3254 756
rect 3080 737 3142 746
rect 3080 703 3100 737
rect 3134 703 3142 737
rect 3080 694 3142 703
rect 3194 737 3254 746
rect 3194 703 3208 737
rect 3242 703 3254 737
rect 3194 694 3254 703
rect 3080 684 3254 694
rect 3656 746 3830 756
rect 3656 737 3718 746
rect 3656 703 3676 737
rect 3710 703 3718 737
rect 3656 694 3718 703
rect 3770 737 3830 746
rect 3770 703 3784 737
rect 3818 703 3830 737
rect 3770 694 3830 703
rect 3656 684 3830 694
rect 4232 746 4406 756
rect 4232 737 4294 746
rect 4232 703 4252 737
rect 4286 703 4294 737
rect 4232 694 4294 703
rect 4346 737 4406 746
rect 4346 703 4360 737
rect 4394 703 4406 737
rect 4346 694 4406 703
rect 4232 684 4406 694
rect 5960 746 6134 756
rect 5960 737 6022 746
rect 5960 703 5980 737
rect 6014 703 6022 737
rect 5960 694 6022 703
rect 6074 737 6134 746
rect 6074 703 6088 737
rect 6122 703 6134 737
rect 6074 694 6134 703
rect 5960 684 6134 694
rect 6536 746 6710 756
rect 6536 737 6598 746
rect 6536 703 6556 737
rect 6590 703 6598 737
rect 6536 694 6598 703
rect 6650 737 6710 746
rect 6650 703 6664 737
rect 6698 703 6710 737
rect 6650 694 6710 703
rect 6536 684 6710 694
rect 7112 746 7286 756
rect 7112 737 7174 746
rect 7112 703 7132 737
rect 7166 703 7174 737
rect 7112 694 7174 703
rect 7226 737 7286 746
rect 7226 703 7240 737
rect 7274 703 7286 737
rect 7226 694 7286 703
rect 7112 684 7286 694
rect 7688 746 7862 756
rect 7688 737 7750 746
rect 7688 703 7708 737
rect 7742 703 7750 737
rect 7688 694 7750 703
rect 7802 737 7862 746
rect 7802 703 7816 737
rect 7850 703 7862 737
rect 7802 694 7862 703
rect 7688 684 7862 694
rect 8174 738 8264 756
rect 8174 702 8196 738
rect 8232 702 8264 738
rect 8174 684 8264 702
rect 8438 746 8528 756
rect 8438 694 8470 746
rect 8522 694 8528 746
rect 8438 684 8528 694
rect 9416 746 9590 756
rect 9416 737 9478 746
rect 9416 703 9436 737
rect 9470 703 9478 737
rect 9416 694 9478 703
rect 9530 737 9590 746
rect 9530 703 9544 737
rect 9578 703 9590 737
rect 9530 694 9590 703
rect 9416 684 9590 694
rect 9992 746 10166 756
rect 9992 737 10054 746
rect 9992 703 10012 737
rect 10046 703 10054 737
rect 9992 694 10054 703
rect 10106 737 10166 746
rect 10106 703 10120 737
rect 10154 703 10166 737
rect 10106 694 10166 703
rect 9992 684 10166 694
rect 10568 746 10742 756
rect 10568 737 10630 746
rect 10568 703 10588 737
rect 10622 703 10630 737
rect 10568 694 10630 703
rect 10682 737 10742 746
rect 10682 703 10696 737
rect 10730 703 10742 737
rect 10682 694 10742 703
rect 10568 684 10742 694
rect 11054 738 11144 756
rect 11054 702 11076 738
rect 11112 702 11144 738
rect 11054 684 11144 702
rect 11318 746 11408 756
rect 11318 694 11350 746
rect 11402 694 11408 746
rect 11318 684 11408 694
rect 12008 746 12182 756
rect 12008 737 12070 746
rect 12008 703 12028 737
rect 12062 703 12070 737
rect 12008 694 12070 703
rect 12122 737 12182 746
rect 12122 703 12136 737
rect 12170 703 12182 737
rect 12122 694 12182 703
rect 12008 684 12182 694
rect 12584 746 12758 756
rect 12584 737 12646 746
rect 12584 703 12604 737
rect 12638 703 12646 737
rect 12584 694 12646 703
rect 12698 737 12758 746
rect 12698 703 12712 737
rect 12746 703 12758 737
rect 12698 694 12758 703
rect 12584 684 12758 694
rect 13160 746 13334 756
rect 13160 737 13222 746
rect 13160 703 13180 737
rect 13214 703 13222 737
rect 13160 694 13222 703
rect 13274 737 13334 746
rect 13274 703 13288 737
rect 13322 703 13334 737
rect 13274 694 13334 703
rect 13160 684 13334 694
rect 13736 746 13910 756
rect 13736 737 13798 746
rect 13736 703 13756 737
rect 13790 703 13798 737
rect 13736 694 13798 703
rect 13850 737 13910 746
rect 13850 703 13864 737
rect 13898 703 13910 737
rect 13850 694 13910 703
rect 13736 684 13910 694
rect 14888 746 15062 756
rect 14888 737 14950 746
rect 14888 703 14908 737
rect 14942 703 14950 737
rect 14888 694 14950 703
rect 15002 737 15062 746
rect 15002 703 15016 737
rect 15050 703 15062 737
rect 15002 694 15062 703
rect 14888 684 15062 694
rect 15466 746 15640 756
rect 15466 737 15526 746
rect 15466 703 15478 737
rect 15512 703 15526 737
rect 15466 694 15526 703
rect 15578 737 15640 746
rect 15578 703 15586 737
rect 15620 703 15640 737
rect 15578 694 15640 703
rect 15466 684 15640 694
rect 16040 746 16214 756
rect 16040 737 16102 746
rect 16040 703 16060 737
rect 16094 703 16102 737
rect 16040 694 16102 703
rect 16154 737 16214 746
rect 16154 703 16168 737
rect 16202 703 16214 737
rect 16154 694 16214 703
rect 16040 684 16214 694
rect 16328 746 16502 756
rect 16328 737 16390 746
rect 16328 703 16348 737
rect 16382 703 16390 737
rect 16328 694 16390 703
rect 16442 737 16502 746
rect 16442 703 16456 737
rect 16490 703 16502 737
rect 16442 694 16502 703
rect 16328 684 16502 694
rect 17480 746 17654 756
rect 17480 737 17542 746
rect 17480 703 17500 737
rect 17534 703 17542 737
rect 17480 694 17542 703
rect 17594 737 17654 746
rect 17594 703 17608 737
rect 17642 703 17654 737
rect 17594 694 17654 703
rect 17480 684 17654 694
rect 17768 746 17942 756
rect 17768 737 17830 746
rect 17768 703 17788 737
rect 17822 703 17830 737
rect 17768 694 17830 703
rect 17882 737 17942 746
rect 17882 703 17896 737
rect 17930 703 17942 737
rect 17882 694 17942 703
rect 17768 684 17942 694
rect 18056 746 18230 756
rect 18056 737 18118 746
rect 18056 703 18076 737
rect 18110 703 18118 737
rect 18056 694 18118 703
rect 18170 737 18230 746
rect 18170 703 18184 737
rect 18218 703 18230 737
rect 18170 694 18230 703
rect 18056 684 18230 694
rect 18344 746 18518 756
rect 18344 737 18406 746
rect 18344 703 18364 737
rect 18398 703 18406 737
rect 18344 694 18406 703
rect 18458 737 18518 746
rect 18458 703 18472 737
rect 18506 703 18518 737
rect 18458 694 18518 703
rect 18344 684 18518 694
rect 18632 746 18806 756
rect 18632 737 18694 746
rect 18632 703 18652 737
rect 18686 703 18694 737
rect 18632 694 18694 703
rect 18746 737 18806 746
rect 18746 703 18760 737
rect 18794 703 18806 737
rect 18746 694 18806 703
rect 18632 684 18806 694
rect 18920 746 19094 756
rect 18920 737 18982 746
rect 18920 703 18940 737
rect 18974 703 18982 737
rect 18920 694 18982 703
rect 19034 737 19094 746
rect 19034 703 19048 737
rect 19082 703 19094 737
rect 19034 694 19094 703
rect 18920 684 19094 694
rect 19208 746 19382 756
rect 19208 737 19270 746
rect 19208 703 19228 737
rect 19262 703 19270 737
rect 19208 694 19270 703
rect 19322 737 19382 746
rect 19322 703 19336 737
rect 19370 703 19382 737
rect 19322 694 19382 703
rect 19208 684 19382 694
rect 19496 746 19670 756
rect 19496 737 19558 746
rect 19496 703 19516 737
rect 19550 703 19558 737
rect 19496 694 19558 703
rect 19610 737 19670 746
rect 19610 703 19624 737
rect 19658 703 19670 737
rect 19610 694 19670 703
rect 19496 684 19670 694
rect 19784 746 19958 756
rect 19784 737 19846 746
rect 19784 703 19804 737
rect 19838 703 19846 737
rect 19784 694 19846 703
rect 19898 737 19958 746
rect 19898 703 19912 737
rect 19946 703 19958 737
rect 19898 694 19958 703
rect 19784 684 19958 694
rect 20072 746 20246 756
rect 20072 737 20134 746
rect 20072 703 20092 737
rect 20126 703 20134 737
rect 20072 694 20134 703
rect 20186 737 20246 746
rect 20186 703 20200 737
rect 20234 703 20246 737
rect 20186 694 20246 703
rect 20072 684 20246 694
rect 20360 746 20534 756
rect 20360 737 20422 746
rect 20360 703 20380 737
rect 20414 703 20422 737
rect 20360 694 20422 703
rect 20474 737 20534 746
rect 20474 703 20488 737
rect 20522 703 20534 737
rect 20474 694 20534 703
rect 20360 684 20534 694
rect 20648 746 20822 756
rect 20648 737 20710 746
rect 20648 703 20668 737
rect 20702 703 20710 737
rect 20648 694 20710 703
rect 20762 737 20822 746
rect 20762 703 20776 737
rect 20810 703 20822 737
rect 20762 694 20822 703
rect 20648 684 20822 694
rect 690 578 750 594
rect 690 538 700 578
rect 740 538 750 578
rect 114 480 174 504
rect 114 328 124 480
rect 164 328 174 480
rect 258 480 318 504
rect 258 464 268 480
rect 256 458 268 464
rect 308 464 318 480
rect 402 480 462 504
rect 308 458 320 464
rect 256 406 262 458
rect 314 406 320 458
rect 256 400 268 406
rect 114 32 174 328
rect 258 328 268 400
rect 308 400 320 406
rect 308 328 318 400
rect 258 188 318 328
rect 402 328 412 480
rect 452 328 462 480
rect 402 32 462 328
rect 690 478 750 538
rect 690 438 700 478
rect 740 438 750 478
rect 834 578 894 594
rect 834 538 844 578
rect 884 538 894 578
rect 834 478 894 538
rect 834 464 844 478
rect 690 378 750 438
rect 832 458 844 464
rect 884 464 894 478
rect 978 578 1038 594
rect 978 538 988 578
rect 1028 538 1038 578
rect 978 478 1038 538
rect 884 458 896 464
rect 832 406 838 458
rect 890 406 896 458
rect 832 400 896 406
rect 978 438 988 478
rect 1028 438 1038 478
rect 690 338 700 378
rect 740 338 750 378
rect 690 278 750 338
rect 690 238 700 278
rect 740 238 750 278
rect 690 32 750 238
rect 834 378 894 400
rect 834 338 844 378
rect 884 338 894 378
rect 834 278 894 338
rect 834 238 844 278
rect 884 238 894 278
rect 834 188 894 238
rect 978 378 1038 438
rect 978 338 988 378
rect 1028 338 1038 378
rect 978 278 1038 338
rect 978 238 988 278
rect 1028 238 1038 278
rect 978 32 1038 238
rect 1266 578 1326 594
rect 1266 538 1276 578
rect 1316 538 1326 578
rect 1266 478 1326 538
rect 1266 438 1276 478
rect 1316 438 1326 478
rect 1410 578 1470 594
rect 1410 538 1420 578
rect 1460 538 1470 578
rect 1410 478 1470 538
rect 1410 464 1420 478
rect 1266 378 1326 438
rect 1408 458 1420 464
rect 1460 464 1470 478
rect 1554 578 1614 594
rect 1554 538 1564 578
rect 1604 538 1614 578
rect 1554 478 1614 538
rect 1460 458 1472 464
rect 1408 406 1414 458
rect 1466 406 1472 458
rect 1408 400 1472 406
rect 1554 438 1564 478
rect 1604 438 1614 478
rect 1266 338 1276 378
rect 1316 338 1326 378
rect 1266 278 1326 338
rect 1266 238 1276 278
rect 1316 238 1326 278
rect 1266 32 1326 238
rect 1410 378 1470 400
rect 1410 338 1420 378
rect 1460 338 1470 378
rect 1410 278 1470 338
rect 1410 238 1420 278
rect 1460 238 1470 278
rect 1410 188 1470 238
rect 1554 378 1614 438
rect 1554 338 1564 378
rect 1604 338 1614 378
rect 1554 278 1614 338
rect 1842 578 1902 594
rect 1842 538 1852 578
rect 1892 538 1902 578
rect 1842 478 1902 538
rect 1842 438 1852 478
rect 1892 438 1902 478
rect 1986 578 2046 594
rect 1986 538 1996 578
rect 2036 538 2046 578
rect 1986 478 2046 538
rect 1986 464 1996 478
rect 1842 378 1902 438
rect 1984 458 1996 464
rect 2036 464 2046 478
rect 2130 578 2190 594
rect 2130 538 2140 578
rect 2180 538 2190 578
rect 2130 478 2190 538
rect 2036 458 2048 464
rect 1984 406 1990 458
rect 2042 406 2048 458
rect 1984 400 2048 406
rect 2130 438 2140 478
rect 2180 438 2190 478
rect 1842 338 1852 378
rect 1892 338 1902 378
rect 1842 320 1902 338
rect 1986 378 2046 400
rect 1986 338 1996 378
rect 2036 338 2046 378
rect 1554 238 1564 278
rect 1604 238 1614 278
rect 1840 314 1904 320
rect 1840 262 1846 314
rect 1898 262 1904 314
rect 1840 256 1852 262
rect 1554 32 1614 238
rect 1842 238 1852 256
rect 1892 256 1904 262
rect 1986 278 2046 338
rect 2130 378 2190 438
rect 2130 338 2140 378
rect 2180 338 2190 378
rect 2130 320 2190 338
rect 2994 578 3054 594
rect 2994 538 3004 578
rect 3044 538 3054 578
rect 2994 478 3054 538
rect 2994 438 3004 478
rect 3044 438 3054 478
rect 3138 578 3198 594
rect 3138 538 3148 578
rect 3188 538 3198 578
rect 3138 478 3198 538
rect 3138 464 3148 478
rect 2994 378 3054 438
rect 3136 458 3148 464
rect 3188 464 3198 478
rect 3282 578 3342 594
rect 3282 538 3292 578
rect 3332 538 3342 578
rect 3282 478 3342 538
rect 3188 458 3200 464
rect 3136 406 3142 458
rect 3194 406 3200 458
rect 3136 400 3200 406
rect 3282 438 3292 478
rect 3332 438 3342 478
rect 2994 338 3004 378
rect 3044 338 3054 378
rect 2994 320 3054 338
rect 3138 378 3198 400
rect 3138 338 3148 378
rect 3188 338 3198 378
rect 1892 238 1902 256
rect 1842 188 1902 238
rect 1986 238 1996 278
rect 2036 238 2046 278
rect 2128 314 2192 320
rect 2128 262 2134 314
rect 2186 262 2192 314
rect 2128 256 2140 262
rect 1986 188 2046 238
rect 2130 238 2140 256
rect 2180 256 2192 262
rect 2992 314 3056 320
rect 2992 262 2998 314
rect 3050 262 3056 314
rect 2992 256 3004 262
rect 2180 238 2190 256
rect 2130 188 2190 238
rect 2994 238 3004 256
rect 3044 256 3056 262
rect 3138 278 3198 338
rect 3282 378 3342 438
rect 3282 338 3292 378
rect 3332 338 3342 378
rect 3282 320 3342 338
rect 3570 578 3630 594
rect 3570 538 3580 578
rect 3620 538 3630 578
rect 3570 478 3630 538
rect 3570 438 3580 478
rect 3620 438 3630 478
rect 3714 578 3774 594
rect 3714 538 3724 578
rect 3764 538 3774 578
rect 3714 478 3774 538
rect 3714 464 3724 478
rect 3570 378 3630 438
rect 3712 458 3724 464
rect 3764 464 3774 478
rect 3858 578 3918 594
rect 3858 538 3868 578
rect 3908 538 3918 578
rect 3858 478 3918 538
rect 3764 458 3776 464
rect 3712 406 3718 458
rect 3770 406 3776 458
rect 3712 400 3776 406
rect 3858 438 3868 478
rect 3908 438 3918 478
rect 3570 338 3580 378
rect 3620 338 3630 378
rect 3044 238 3054 256
rect 2994 188 3054 238
rect 3138 238 3148 278
rect 3188 238 3198 278
rect 3280 314 3344 320
rect 3280 262 3286 314
rect 3338 262 3344 314
rect 3280 256 3292 262
rect 3138 188 3198 238
rect 3282 238 3292 256
rect 3332 256 3344 262
rect 3570 278 3630 338
rect 3332 238 3342 256
rect 3282 188 3342 238
rect 3570 238 3580 278
rect 3620 238 3630 278
rect 3570 32 3630 238
rect 3714 378 3774 400
rect 3714 338 3724 378
rect 3764 338 3774 378
rect 3714 278 3774 338
rect 3714 238 3724 278
rect 3764 238 3774 278
rect 3714 188 3774 238
rect 3858 378 3918 438
rect 3858 338 3868 378
rect 3908 338 3918 378
rect 3858 278 3918 338
rect 3858 238 3868 278
rect 3908 238 3918 278
rect 3858 32 3918 238
rect 4146 578 4206 594
rect 4146 538 4156 578
rect 4196 538 4206 578
rect 4146 478 4206 538
rect 4146 438 4156 478
rect 4196 438 4206 478
rect 4290 578 4350 594
rect 4290 538 4300 578
rect 4340 538 4350 578
rect 4290 478 4350 538
rect 4290 464 4300 478
rect 4146 378 4206 438
rect 4288 458 4300 464
rect 4340 464 4350 478
rect 4434 578 4494 594
rect 4434 538 4444 578
rect 4484 538 4494 578
rect 4434 478 4494 538
rect 5874 578 5934 594
rect 5874 538 5884 578
rect 5924 538 5934 578
rect 4340 458 4352 464
rect 4288 406 4294 458
rect 4346 406 4352 458
rect 4288 400 4352 406
rect 4434 438 4444 478
rect 4484 438 4494 478
rect 4146 338 4156 378
rect 4196 338 4206 378
rect 4146 278 4206 338
rect 4146 238 4156 278
rect 4196 238 4206 278
rect 4146 32 4206 238
rect 4290 378 4350 400
rect 4290 338 4300 378
rect 4340 338 4350 378
rect 4290 278 4350 338
rect 4290 238 4300 278
rect 4340 238 4350 278
rect 4290 188 4350 238
rect 4434 378 4494 438
rect 4434 338 4444 378
rect 4484 338 4494 378
rect 4434 278 4494 338
rect 4434 238 4444 278
rect 4484 238 4494 278
rect 4434 32 4494 238
rect 4722 480 4782 504
rect 4722 328 4732 480
rect 4772 328 4782 480
rect 4866 480 4926 504
rect 4866 464 4876 480
rect 4864 458 4876 464
rect 4916 464 4926 480
rect 5010 480 5070 504
rect 4916 458 4928 464
rect 4864 406 4870 458
rect 4922 406 4928 458
rect 4864 400 4876 406
rect 4722 32 4782 328
rect 4866 328 4876 400
rect 4916 400 4928 406
rect 4916 328 4926 400
rect 4866 188 4926 328
rect 5010 328 5020 480
rect 5060 328 5070 480
rect 5010 32 5070 328
rect 5298 480 5358 504
rect 5298 328 5308 480
rect 5348 328 5358 480
rect 5442 480 5502 504
rect 5442 464 5452 480
rect 5440 458 5452 464
rect 5492 464 5502 480
rect 5586 480 5646 504
rect 5492 458 5504 464
rect 5440 406 5446 458
rect 5498 406 5504 458
rect 5440 400 5452 406
rect 5298 32 5358 328
rect 5442 328 5452 400
rect 5492 400 5504 406
rect 5492 328 5502 400
rect 5442 188 5502 328
rect 5586 328 5596 480
rect 5636 328 5646 480
rect 5586 32 5646 328
rect 5874 478 5934 538
rect 5874 438 5884 478
rect 5924 438 5934 478
rect 6018 578 6078 594
rect 6018 538 6028 578
rect 6068 538 6078 578
rect 6018 478 6078 538
rect 6018 464 6028 478
rect 5874 378 5934 438
rect 6016 458 6028 464
rect 6068 464 6078 478
rect 6162 578 6222 594
rect 6162 538 6172 578
rect 6212 538 6222 578
rect 6162 478 6222 538
rect 6068 458 6080 464
rect 6016 406 6022 458
rect 6074 406 6080 458
rect 6016 400 6080 406
rect 6162 438 6172 478
rect 6212 438 6222 478
rect 5874 338 5884 378
rect 5924 338 5934 378
rect 5874 278 5934 338
rect 5874 238 5884 278
rect 5924 238 5934 278
rect 5874 32 5934 238
rect 6018 378 6078 400
rect 6018 338 6028 378
rect 6068 338 6078 378
rect 6018 278 6078 338
rect 6018 238 6028 278
rect 6068 238 6078 278
rect 6018 188 6078 238
rect 6162 378 6222 438
rect 6162 338 6172 378
rect 6212 338 6222 378
rect 6162 278 6222 338
rect 6162 238 6172 278
rect 6212 238 6222 278
rect 6162 32 6222 238
rect 6450 578 6510 594
rect 6450 538 6460 578
rect 6500 538 6510 578
rect 6450 478 6510 538
rect 6450 438 6460 478
rect 6500 438 6510 478
rect 6594 578 6654 594
rect 6594 538 6604 578
rect 6644 538 6654 578
rect 6594 478 6654 538
rect 6594 464 6604 478
rect 6450 378 6510 438
rect 6592 458 6604 464
rect 6644 464 6654 478
rect 6738 578 6798 594
rect 6738 538 6748 578
rect 6788 538 6798 578
rect 6738 478 6798 538
rect 6644 458 6656 464
rect 6592 406 6598 458
rect 6650 406 6656 458
rect 6592 400 6656 406
rect 6738 438 6748 478
rect 6788 438 6798 478
rect 6450 338 6460 378
rect 6500 338 6510 378
rect 6450 278 6510 338
rect 6450 238 6460 278
rect 6500 238 6510 278
rect 6450 32 6510 238
rect 6594 378 6654 400
rect 6594 338 6604 378
rect 6644 338 6654 378
rect 6594 278 6654 338
rect 6594 238 6604 278
rect 6644 238 6654 278
rect 6594 188 6654 238
rect 6738 378 6798 438
rect 6738 338 6748 378
rect 6788 338 6798 378
rect 6738 278 6798 338
rect 6738 238 6748 278
rect 6788 238 6798 278
rect 6738 32 6798 238
rect 7026 578 7086 594
rect 7026 538 7036 578
rect 7076 538 7086 578
rect 7026 478 7086 538
rect 7026 438 7036 478
rect 7076 438 7086 478
rect 7170 578 7230 594
rect 7170 538 7180 578
rect 7220 538 7230 578
rect 7170 478 7230 538
rect 7170 464 7180 478
rect 7026 378 7086 438
rect 7168 458 7180 464
rect 7220 464 7230 478
rect 7314 578 7374 594
rect 7314 538 7324 578
rect 7364 538 7374 578
rect 7314 478 7374 538
rect 7220 458 7232 464
rect 7168 406 7174 458
rect 7226 406 7232 458
rect 7168 400 7232 406
rect 7314 438 7324 478
rect 7364 438 7374 478
rect 7602 578 7662 594
rect 7602 538 7612 578
rect 7652 538 7662 578
rect 7602 478 7662 538
rect 7602 464 7612 478
rect 7026 338 7036 378
rect 7076 338 7086 378
rect 7026 278 7086 338
rect 7026 238 7036 278
rect 7076 238 7086 278
rect 7026 32 7086 238
rect 7170 378 7230 400
rect 7170 338 7180 378
rect 7220 338 7230 378
rect 7170 278 7230 338
rect 7170 238 7180 278
rect 7220 238 7230 278
rect 7170 188 7230 238
rect 7314 378 7374 438
rect 7600 458 7612 464
rect 7652 464 7662 478
rect 7746 578 7806 594
rect 7746 538 7756 578
rect 7796 538 7806 578
rect 7746 478 7806 538
rect 7652 458 7664 464
rect 7600 406 7606 458
rect 7658 406 7664 458
rect 7600 400 7664 406
rect 7746 438 7756 478
rect 7796 438 7806 478
rect 7890 578 7950 594
rect 7890 538 7900 578
rect 7940 538 7950 578
rect 7890 478 7950 538
rect 7890 464 7900 478
rect 7314 338 7324 378
rect 7364 338 7374 378
rect 7314 278 7374 338
rect 7314 238 7324 278
rect 7364 238 7374 278
rect 7314 32 7374 238
rect 7602 378 7662 400
rect 7602 338 7612 378
rect 7652 338 7662 378
rect 7602 278 7662 338
rect 7746 378 7806 438
rect 7888 458 7900 464
rect 7940 464 7950 478
rect 8178 578 8238 594
rect 8178 538 8188 578
rect 8228 538 8238 578
rect 8178 478 8238 538
rect 7940 458 7952 464
rect 7888 406 7894 458
rect 7946 406 7952 458
rect 7888 400 7952 406
rect 8178 438 8188 478
rect 8228 438 8238 478
rect 7746 338 7756 378
rect 7796 338 7806 378
rect 7746 320 7806 338
rect 7890 378 7950 400
rect 7890 338 7900 378
rect 7940 338 7950 378
rect 7602 238 7612 278
rect 7652 238 7662 278
rect 7744 314 7808 320
rect 7744 262 7750 314
rect 7802 262 7808 314
rect 7744 256 7756 262
rect 7602 188 7662 238
rect 7746 238 7756 256
rect 7796 256 7808 262
rect 7890 278 7950 338
rect 7796 238 7806 256
rect 7746 188 7806 238
rect 7890 238 7900 278
rect 7940 238 7950 278
rect 7890 188 7950 238
rect 8178 378 8238 438
rect 8178 338 8188 378
rect 8228 338 8238 378
rect 8178 278 8238 338
rect 8178 238 8188 278
rect 8228 238 8238 278
rect 8178 32 8238 238
rect 8322 578 8382 594
rect 8322 538 8332 578
rect 8372 538 8382 578
rect 8322 478 8382 538
rect 8322 438 8332 478
rect 8372 438 8382 478
rect 8322 378 8382 438
rect 8322 338 8332 378
rect 8372 338 8382 378
rect 8322 278 8382 338
rect 8466 578 8526 594
rect 8466 538 8476 578
rect 8516 538 8526 578
rect 8466 478 8526 538
rect 9330 578 9390 594
rect 9330 538 9340 578
rect 9380 538 9390 578
rect 8466 438 8476 478
rect 8516 438 8526 478
rect 8466 378 8526 438
rect 8466 338 8476 378
rect 8516 338 8526 378
rect 8466 320 8526 338
rect 8754 480 8814 504
rect 8754 328 8764 480
rect 8804 328 8814 480
rect 8898 480 8958 504
rect 8898 464 8908 480
rect 8896 458 8908 464
rect 8948 464 8958 480
rect 9042 480 9102 504
rect 8948 458 8960 464
rect 8896 406 8902 458
rect 8954 406 8960 458
rect 8896 400 8908 406
rect 8322 238 8332 278
rect 8372 238 8382 278
rect 8464 314 8528 320
rect 8464 262 8470 314
rect 8522 262 8528 314
rect 8464 256 8476 262
rect 8322 188 8382 238
rect 8466 238 8476 256
rect 8516 256 8528 262
rect 8516 238 8526 256
rect 8466 188 8526 238
rect 8754 32 8814 328
rect 8898 328 8908 400
rect 8948 400 8960 406
rect 8948 328 8958 400
rect 8898 188 8958 328
rect 9042 328 9052 480
rect 9092 328 9102 480
rect 9042 32 9102 328
rect 9330 478 9390 538
rect 9330 438 9340 478
rect 9380 438 9390 478
rect 9474 578 9534 594
rect 9474 538 9484 578
rect 9524 538 9534 578
rect 9474 478 9534 538
rect 9474 464 9484 478
rect 9330 378 9390 438
rect 9472 458 9484 464
rect 9524 464 9534 478
rect 9618 578 9678 594
rect 9618 538 9628 578
rect 9668 538 9678 578
rect 9618 478 9678 538
rect 9524 458 9536 464
rect 9472 406 9478 458
rect 9530 406 9536 458
rect 9472 400 9536 406
rect 9618 438 9628 478
rect 9668 438 9678 478
rect 9330 338 9340 378
rect 9380 338 9390 378
rect 9330 278 9390 338
rect 9330 238 9340 278
rect 9380 238 9390 278
rect 9330 32 9390 238
rect 9474 378 9534 400
rect 9474 338 9484 378
rect 9524 338 9534 378
rect 9474 278 9534 338
rect 9474 238 9484 278
rect 9524 238 9534 278
rect 9474 188 9534 238
rect 9618 378 9678 438
rect 9618 338 9628 378
rect 9668 338 9678 378
rect 9618 278 9678 338
rect 9618 238 9628 278
rect 9668 238 9678 278
rect 9618 32 9678 238
rect 9906 578 9966 594
rect 9906 538 9916 578
rect 9956 538 9966 578
rect 9906 478 9966 538
rect 9906 438 9916 478
rect 9956 438 9966 478
rect 10050 578 10110 594
rect 10050 538 10060 578
rect 10100 538 10110 578
rect 10050 478 10110 538
rect 10050 464 10060 478
rect 9906 378 9966 438
rect 10048 458 10060 464
rect 10100 464 10110 478
rect 10194 578 10254 594
rect 10194 538 10204 578
rect 10244 538 10254 578
rect 10194 478 10254 538
rect 10100 458 10112 464
rect 10048 406 10054 458
rect 10106 406 10112 458
rect 10048 400 10112 406
rect 10194 438 10204 478
rect 10244 438 10254 478
rect 10482 578 10542 594
rect 10482 538 10492 578
rect 10532 538 10542 578
rect 10482 478 10542 538
rect 10482 464 10492 478
rect 9906 338 9916 378
rect 9956 338 9966 378
rect 9906 278 9966 338
rect 9906 238 9916 278
rect 9956 238 9966 278
rect 9906 32 9966 238
rect 10050 378 10110 400
rect 10050 338 10060 378
rect 10100 338 10110 378
rect 10050 278 10110 338
rect 10050 238 10060 278
rect 10100 238 10110 278
rect 10050 188 10110 238
rect 10194 378 10254 438
rect 10480 458 10492 464
rect 10532 464 10542 478
rect 10626 578 10686 594
rect 10626 538 10636 578
rect 10676 538 10686 578
rect 10626 478 10686 538
rect 10532 458 10544 464
rect 10480 406 10486 458
rect 10538 406 10544 458
rect 10480 400 10544 406
rect 10626 438 10636 478
rect 10676 438 10686 478
rect 10770 578 10830 594
rect 10770 538 10780 578
rect 10820 538 10830 578
rect 10770 478 10830 538
rect 10770 464 10780 478
rect 10194 338 10204 378
rect 10244 338 10254 378
rect 10194 278 10254 338
rect 10194 238 10204 278
rect 10244 238 10254 278
rect 10194 32 10254 238
rect 10482 378 10542 400
rect 10482 338 10492 378
rect 10532 338 10542 378
rect 10482 278 10542 338
rect 10626 378 10686 438
rect 10768 458 10780 464
rect 10820 464 10830 478
rect 11058 578 11118 594
rect 11058 538 11068 578
rect 11108 538 11118 578
rect 11058 478 11118 538
rect 10820 458 10832 464
rect 10768 406 10774 458
rect 10826 406 10832 458
rect 10768 400 10832 406
rect 11058 438 11068 478
rect 11108 438 11118 478
rect 10626 338 10636 378
rect 10676 338 10686 378
rect 10626 320 10686 338
rect 10770 378 10830 400
rect 10770 338 10780 378
rect 10820 338 10830 378
rect 10482 238 10492 278
rect 10532 238 10542 278
rect 10624 314 10688 320
rect 10624 262 10630 314
rect 10682 262 10688 314
rect 10624 256 10636 262
rect 10482 188 10542 238
rect 10626 238 10636 256
rect 10676 256 10688 262
rect 10770 278 10830 338
rect 10676 238 10686 256
rect 10626 188 10686 238
rect 10770 238 10780 278
rect 10820 238 10830 278
rect 10770 188 10830 238
rect 11058 378 11118 438
rect 11058 338 11068 378
rect 11108 338 11118 378
rect 11058 278 11118 338
rect 11058 238 11068 278
rect 11108 238 11118 278
rect 11058 32 11118 238
rect 11202 578 11262 594
rect 11202 538 11212 578
rect 11252 538 11262 578
rect 11202 478 11262 538
rect 11202 438 11212 478
rect 11252 438 11262 478
rect 11202 378 11262 438
rect 11202 338 11212 378
rect 11252 338 11262 378
rect 11202 278 11262 338
rect 11346 578 11406 594
rect 11346 538 11356 578
rect 11396 538 11406 578
rect 11346 478 11406 538
rect 11346 438 11356 478
rect 11396 438 11406 478
rect 11346 378 11406 438
rect 11346 338 11356 378
rect 11396 338 11406 378
rect 11346 320 11406 338
rect 11922 578 11982 594
rect 11922 538 11932 578
rect 11972 538 11982 578
rect 11922 478 11982 538
rect 11922 438 11932 478
rect 11972 438 11982 478
rect 12066 578 12126 594
rect 12066 538 12076 578
rect 12116 538 12126 578
rect 12066 478 12126 538
rect 12066 464 12076 478
rect 11922 378 11982 438
rect 12064 458 12076 464
rect 12116 464 12126 478
rect 12210 578 12270 594
rect 12210 538 12220 578
rect 12260 538 12270 578
rect 12210 478 12270 538
rect 12116 458 12128 464
rect 12064 406 12070 458
rect 12122 406 12128 458
rect 12064 400 12128 406
rect 12210 438 12220 478
rect 12260 438 12270 478
rect 11922 338 11932 378
rect 11972 338 11982 378
rect 11202 238 11212 278
rect 11252 238 11262 278
rect 11344 314 11408 320
rect 11344 262 11350 314
rect 11402 262 11408 314
rect 11344 256 11356 262
rect 11202 188 11262 238
rect 11346 238 11356 256
rect 11396 256 11408 262
rect 11922 278 11982 338
rect 11396 238 11406 256
rect 11346 188 11406 238
rect 11922 238 11932 278
rect 11972 238 11982 278
rect 11922 32 11982 238
rect 12066 378 12126 400
rect 12066 338 12076 378
rect 12116 338 12126 378
rect 12066 278 12126 338
rect 12066 238 12076 278
rect 12116 238 12126 278
rect 12066 188 12126 238
rect 12210 378 12270 438
rect 12210 338 12220 378
rect 12260 338 12270 378
rect 12210 278 12270 338
rect 12210 238 12220 278
rect 12260 238 12270 278
rect 12210 32 12270 238
rect 12498 578 12558 594
rect 12498 538 12508 578
rect 12548 538 12558 578
rect 12498 478 12558 538
rect 12498 438 12508 478
rect 12548 438 12558 478
rect 12642 578 12702 594
rect 12642 538 12652 578
rect 12692 538 12702 578
rect 12642 478 12702 538
rect 12642 464 12652 478
rect 12498 378 12558 438
rect 12640 458 12652 464
rect 12692 464 12702 478
rect 12786 578 12846 594
rect 12786 538 12796 578
rect 12836 538 12846 578
rect 12786 478 12846 538
rect 12692 458 12704 464
rect 12640 406 12646 458
rect 12698 406 12704 458
rect 12640 400 12704 406
rect 12786 438 12796 478
rect 12836 438 12846 478
rect 12498 338 12508 378
rect 12548 338 12558 378
rect 12498 278 12558 338
rect 12498 238 12508 278
rect 12548 238 12558 278
rect 12498 32 12558 238
rect 12642 378 12702 400
rect 12642 338 12652 378
rect 12692 338 12702 378
rect 12642 278 12702 338
rect 12642 238 12652 278
rect 12692 238 12702 278
rect 12642 188 12702 238
rect 12786 378 12846 438
rect 12786 338 12796 378
rect 12836 338 12846 378
rect 12786 278 12846 338
rect 12786 238 12796 278
rect 12836 238 12846 278
rect 12786 32 12846 238
rect 13074 578 13134 594
rect 13074 538 13084 578
rect 13124 538 13134 578
rect 13074 478 13134 538
rect 13074 438 13084 478
rect 13124 438 13134 478
rect 13218 578 13278 594
rect 13218 538 13228 578
rect 13268 538 13278 578
rect 13218 478 13278 538
rect 13218 464 13228 478
rect 13074 378 13134 438
rect 13216 458 13228 464
rect 13268 464 13278 478
rect 13362 578 13422 594
rect 13362 538 13372 578
rect 13412 538 13422 578
rect 13362 478 13422 538
rect 13268 458 13280 464
rect 13216 406 13222 458
rect 13274 406 13280 458
rect 13216 400 13280 406
rect 13362 438 13372 478
rect 13412 438 13422 478
rect 13074 338 13084 378
rect 13124 338 13134 378
rect 13074 278 13134 338
rect 13074 238 13084 278
rect 13124 238 13134 278
rect 13074 32 13134 238
rect 13218 378 13278 400
rect 13218 338 13228 378
rect 13268 338 13278 378
rect 13218 278 13278 338
rect 13218 238 13228 278
rect 13268 238 13278 278
rect 13218 188 13278 238
rect 13362 378 13422 438
rect 13362 338 13372 378
rect 13412 338 13422 378
rect 13362 278 13422 338
rect 13362 238 13372 278
rect 13412 238 13422 278
rect 13362 32 13422 238
rect 13650 578 13710 594
rect 13650 538 13660 578
rect 13700 538 13710 578
rect 13650 478 13710 538
rect 13650 438 13660 478
rect 13700 438 13710 478
rect 13794 578 13854 594
rect 13794 538 13804 578
rect 13844 538 13854 578
rect 13794 478 13854 538
rect 13794 464 13804 478
rect 13650 378 13710 438
rect 13792 458 13804 464
rect 13844 464 13854 478
rect 13938 578 13998 594
rect 13938 538 13948 578
rect 13988 538 13998 578
rect 13938 478 13998 538
rect 14802 578 14862 594
rect 14802 538 14812 578
rect 14852 538 14862 578
rect 13844 458 13856 464
rect 13792 406 13798 458
rect 13850 406 13856 458
rect 13792 400 13856 406
rect 13938 438 13948 478
rect 13988 438 13998 478
rect 13650 338 13660 378
rect 13700 338 13710 378
rect 13650 278 13710 338
rect 13650 238 13660 278
rect 13700 238 13710 278
rect 13650 32 13710 238
rect 13794 378 13854 400
rect 13794 338 13804 378
rect 13844 338 13854 378
rect 13794 278 13854 338
rect 13794 238 13804 278
rect 13844 238 13854 278
rect 13794 188 13854 238
rect 13938 378 13998 438
rect 13938 338 13948 378
rect 13988 338 13998 378
rect 13938 278 13998 338
rect 13938 238 13948 278
rect 13988 238 13998 278
rect 13938 32 13998 238
rect 14226 480 14286 504
rect 14226 328 14236 480
rect 14276 328 14286 480
rect 14370 480 14430 504
rect 14370 464 14380 480
rect 14368 458 14380 464
rect 14420 464 14430 480
rect 14514 480 14574 504
rect 14420 458 14432 464
rect 14368 406 14374 458
rect 14426 406 14432 458
rect 14368 400 14380 406
rect 14226 32 14286 328
rect 14370 328 14380 400
rect 14420 400 14432 406
rect 14420 328 14430 400
rect 14370 188 14430 328
rect 14514 328 14524 480
rect 14564 328 14574 480
rect 14514 32 14574 328
rect 14802 478 14862 538
rect 14802 438 14812 478
rect 14852 438 14862 478
rect 14946 578 15006 594
rect 14946 538 14956 578
rect 14996 538 15006 578
rect 14946 478 15006 538
rect 14946 464 14956 478
rect 14802 378 14862 438
rect 14944 458 14956 464
rect 14996 464 15006 478
rect 15090 578 15150 594
rect 15090 538 15100 578
rect 15140 538 15150 578
rect 15090 478 15150 538
rect 14996 458 15008 464
rect 14944 406 14950 458
rect 15002 406 15008 458
rect 14944 400 15008 406
rect 15090 438 15100 478
rect 15140 438 15150 478
rect 14802 338 14812 378
rect 14852 338 14862 378
rect 14802 278 14862 338
rect 14802 238 14812 278
rect 14852 238 14862 278
rect 14802 32 14862 238
rect 14946 378 15006 400
rect 14946 338 14956 378
rect 14996 338 15006 378
rect 14946 278 15006 338
rect 14946 238 14956 278
rect 14996 238 15006 278
rect 14946 188 15006 238
rect 15090 378 15150 438
rect 15090 338 15100 378
rect 15140 338 15150 378
rect 15090 278 15150 338
rect 15090 238 15100 278
rect 15140 238 15150 278
rect 15090 32 15150 238
rect 15378 578 15438 594
rect 15378 538 15388 578
rect 15428 538 15438 578
rect 15378 478 15438 538
rect 15378 438 15388 478
rect 15428 438 15438 478
rect 15522 578 15582 594
rect 15522 538 15532 578
rect 15572 538 15582 578
rect 15522 478 15582 538
rect 15522 464 15532 478
rect 15378 378 15438 438
rect 15520 458 15532 464
rect 15572 464 15582 478
rect 15666 578 15726 594
rect 15666 538 15676 578
rect 15716 538 15726 578
rect 15666 478 15726 538
rect 15572 458 15584 464
rect 15520 406 15526 458
rect 15578 406 15584 458
rect 15520 400 15584 406
rect 15666 438 15676 478
rect 15716 438 15726 478
rect 15378 338 15388 378
rect 15428 338 15438 378
rect 15378 278 15438 338
rect 15378 238 15388 278
rect 15428 238 15438 278
rect 15378 32 15438 238
rect 15522 378 15582 400
rect 15522 338 15532 378
rect 15572 338 15582 378
rect 15522 278 15582 338
rect 15522 238 15532 278
rect 15572 238 15582 278
rect 15522 188 15582 238
rect 15666 378 15726 438
rect 15666 338 15676 378
rect 15716 338 15726 378
rect 15666 278 15726 338
rect 15666 238 15676 278
rect 15716 238 15726 278
rect 15666 32 15726 238
rect 15954 578 16014 594
rect 15954 538 15964 578
rect 16004 538 16014 578
rect 15954 478 16014 538
rect 15954 438 15964 478
rect 16004 438 16014 478
rect 16098 578 16158 594
rect 16098 538 16108 578
rect 16148 538 16158 578
rect 16098 478 16158 538
rect 16098 464 16108 478
rect 15954 378 16014 438
rect 16096 458 16108 464
rect 16148 464 16158 478
rect 16242 578 16302 594
rect 16242 538 16252 578
rect 16292 538 16302 578
rect 16242 478 16302 538
rect 16148 458 16160 464
rect 16096 406 16102 458
rect 16154 406 16160 458
rect 16096 400 16160 406
rect 16242 438 16252 478
rect 16292 438 16302 478
rect 16386 578 16446 594
rect 16386 538 16396 578
rect 16436 538 16446 578
rect 16386 478 16446 538
rect 16386 464 16396 478
rect 15954 338 15964 378
rect 16004 338 16014 378
rect 15954 278 16014 338
rect 15954 238 15964 278
rect 16004 238 16014 278
rect 15954 32 16014 238
rect 16098 378 16158 400
rect 16098 338 16108 378
rect 16148 338 16158 378
rect 16098 278 16158 338
rect 16098 238 16108 278
rect 16148 238 16158 278
rect 16098 188 16158 238
rect 16242 378 16302 438
rect 16384 458 16396 464
rect 16436 464 16446 478
rect 16530 578 16590 594
rect 16530 538 16540 578
rect 16580 538 16590 578
rect 16530 478 16590 538
rect 17394 578 17454 594
rect 17394 538 17404 578
rect 17444 538 17454 578
rect 16436 458 16448 464
rect 16384 406 16390 458
rect 16442 406 16448 458
rect 16384 400 16448 406
rect 16530 438 16540 478
rect 16580 438 16590 478
rect 16242 338 16252 378
rect 16292 338 16302 378
rect 16242 278 16302 338
rect 16242 238 16252 278
rect 16292 238 16302 278
rect 16242 32 16302 238
rect 16386 378 16446 400
rect 16386 338 16396 378
rect 16436 338 16446 378
rect 16386 278 16446 338
rect 16386 238 16396 278
rect 16436 238 16446 278
rect 16386 188 16446 238
rect 16530 378 16590 438
rect 16530 338 16540 378
rect 16580 338 16590 378
rect 16530 278 16590 338
rect 16530 238 16540 278
rect 16580 238 16590 278
rect 16530 32 16590 238
rect 16818 480 16878 504
rect 16818 328 16828 480
rect 16868 328 16878 480
rect 16962 480 17022 504
rect 16962 464 16972 480
rect 16960 458 16972 464
rect 17012 464 17022 480
rect 17106 480 17166 504
rect 17012 458 17024 464
rect 16960 406 16966 458
rect 17018 406 17024 458
rect 16960 400 16972 406
rect 16818 32 16878 328
rect 16962 328 16972 400
rect 17012 400 17024 406
rect 17012 328 17022 400
rect 16962 188 17022 328
rect 17106 328 17116 480
rect 17156 328 17166 480
rect 17106 32 17166 328
rect 17394 478 17454 538
rect 17394 438 17404 478
rect 17444 438 17454 478
rect 17538 578 17598 594
rect 17538 538 17548 578
rect 17588 538 17598 578
rect 17538 478 17598 538
rect 17538 464 17548 478
rect 17394 378 17454 438
rect 17536 458 17548 464
rect 17588 464 17598 478
rect 17682 578 17742 594
rect 17682 538 17692 578
rect 17732 538 17742 578
rect 17682 478 17742 538
rect 17588 458 17600 464
rect 17536 406 17542 458
rect 17594 406 17600 458
rect 17536 400 17600 406
rect 17682 438 17692 478
rect 17732 438 17742 478
rect 17826 578 17886 594
rect 17826 538 17836 578
rect 17876 538 17886 578
rect 17826 478 17886 538
rect 17826 464 17836 478
rect 17394 338 17404 378
rect 17444 338 17454 378
rect 17394 278 17454 338
rect 17394 238 17404 278
rect 17444 238 17454 278
rect 17394 32 17454 238
rect 17538 378 17598 400
rect 17538 338 17548 378
rect 17588 338 17598 378
rect 17538 278 17598 338
rect 17538 238 17548 278
rect 17588 238 17598 278
rect 17538 188 17598 238
rect 17682 378 17742 438
rect 17824 458 17836 464
rect 17876 464 17886 478
rect 17970 578 18030 594
rect 17970 538 17980 578
rect 18020 538 18030 578
rect 17970 478 18030 538
rect 17876 458 17888 464
rect 17824 406 17830 458
rect 17882 406 17888 458
rect 17824 400 17888 406
rect 17970 438 17980 478
rect 18020 438 18030 478
rect 18114 578 18174 594
rect 18114 538 18124 578
rect 18164 538 18174 578
rect 18114 478 18174 538
rect 18114 464 18124 478
rect 17682 338 17692 378
rect 17732 338 17742 378
rect 17682 278 17742 338
rect 17682 238 17692 278
rect 17732 238 17742 278
rect 17682 32 17742 238
rect 17826 378 17886 400
rect 17826 338 17836 378
rect 17876 338 17886 378
rect 17826 278 17886 338
rect 17826 238 17836 278
rect 17876 238 17886 278
rect 17826 188 17886 238
rect 17970 378 18030 438
rect 18112 458 18124 464
rect 18164 464 18174 478
rect 18258 578 18318 594
rect 18258 538 18268 578
rect 18308 538 18318 578
rect 18258 478 18318 538
rect 18164 458 18176 464
rect 18112 406 18118 458
rect 18170 406 18176 458
rect 18112 400 18176 406
rect 18258 438 18268 478
rect 18308 438 18318 478
rect 18402 578 18462 594
rect 18402 538 18412 578
rect 18452 538 18462 578
rect 18402 478 18462 538
rect 18402 464 18412 478
rect 17970 338 17980 378
rect 18020 338 18030 378
rect 17970 278 18030 338
rect 17970 238 17980 278
rect 18020 238 18030 278
rect 17970 32 18030 238
rect 18114 378 18174 400
rect 18114 338 18124 378
rect 18164 338 18174 378
rect 18114 278 18174 338
rect 18114 238 18124 278
rect 18164 238 18174 278
rect 18114 188 18174 238
rect 18258 378 18318 438
rect 18400 458 18412 464
rect 18452 464 18462 478
rect 18546 578 18606 594
rect 18546 538 18556 578
rect 18596 538 18606 578
rect 18546 478 18606 538
rect 18452 458 18464 464
rect 18400 406 18406 458
rect 18458 406 18464 458
rect 18400 400 18464 406
rect 18546 438 18556 478
rect 18596 438 18606 478
rect 18690 578 18750 594
rect 18690 538 18700 578
rect 18740 538 18750 578
rect 18690 478 18750 538
rect 18690 464 18700 478
rect 18258 338 18268 378
rect 18308 338 18318 378
rect 18258 278 18318 338
rect 18258 238 18268 278
rect 18308 238 18318 278
rect 18258 32 18318 238
rect 18402 378 18462 400
rect 18402 338 18412 378
rect 18452 338 18462 378
rect 18402 278 18462 338
rect 18402 238 18412 278
rect 18452 238 18462 278
rect 18402 188 18462 238
rect 18546 378 18606 438
rect 18688 458 18700 464
rect 18740 464 18750 478
rect 18834 578 18894 594
rect 18834 538 18844 578
rect 18884 538 18894 578
rect 18834 478 18894 538
rect 18740 458 18752 464
rect 18688 406 18694 458
rect 18746 406 18752 458
rect 18688 400 18752 406
rect 18834 438 18844 478
rect 18884 438 18894 478
rect 18978 578 19038 594
rect 18978 538 18988 578
rect 19028 538 19038 578
rect 18978 478 19038 538
rect 18978 464 18988 478
rect 18546 338 18556 378
rect 18596 338 18606 378
rect 18546 278 18606 338
rect 18546 238 18556 278
rect 18596 238 18606 278
rect 18546 32 18606 238
rect 18690 378 18750 400
rect 18690 338 18700 378
rect 18740 338 18750 378
rect 18690 278 18750 338
rect 18690 238 18700 278
rect 18740 238 18750 278
rect 18690 188 18750 238
rect 18834 378 18894 438
rect 18976 458 18988 464
rect 19028 464 19038 478
rect 19122 578 19182 594
rect 19122 538 19132 578
rect 19172 538 19182 578
rect 19122 478 19182 538
rect 19028 458 19040 464
rect 18976 406 18982 458
rect 19034 406 19040 458
rect 18976 400 19040 406
rect 19122 438 19132 478
rect 19172 438 19182 478
rect 19266 578 19326 594
rect 19266 538 19276 578
rect 19316 538 19326 578
rect 19266 478 19326 538
rect 19266 464 19276 478
rect 18834 338 18844 378
rect 18884 338 18894 378
rect 18834 278 18894 338
rect 18834 238 18844 278
rect 18884 238 18894 278
rect 18834 32 18894 238
rect 18978 378 19038 400
rect 18978 338 18988 378
rect 19028 338 19038 378
rect 18978 278 19038 338
rect 18978 238 18988 278
rect 19028 238 19038 278
rect 18978 188 19038 238
rect 19122 378 19182 438
rect 19264 458 19276 464
rect 19316 464 19326 478
rect 19410 578 19470 594
rect 19410 538 19420 578
rect 19460 538 19470 578
rect 19410 478 19470 538
rect 19316 458 19328 464
rect 19264 406 19270 458
rect 19322 406 19328 458
rect 19264 400 19328 406
rect 19410 438 19420 478
rect 19460 438 19470 478
rect 19554 578 19614 594
rect 19554 538 19564 578
rect 19604 538 19614 578
rect 19554 478 19614 538
rect 19554 464 19564 478
rect 19122 338 19132 378
rect 19172 338 19182 378
rect 19122 278 19182 338
rect 19122 238 19132 278
rect 19172 238 19182 278
rect 19122 32 19182 238
rect 19266 378 19326 400
rect 19266 338 19276 378
rect 19316 338 19326 378
rect 19266 278 19326 338
rect 19266 238 19276 278
rect 19316 238 19326 278
rect 19266 188 19326 238
rect 19410 378 19470 438
rect 19552 458 19564 464
rect 19604 464 19614 478
rect 19698 578 19758 594
rect 19698 538 19708 578
rect 19748 538 19758 578
rect 19698 478 19758 538
rect 19604 458 19616 464
rect 19552 406 19558 458
rect 19610 406 19616 458
rect 19552 400 19616 406
rect 19698 438 19708 478
rect 19748 438 19758 478
rect 19842 578 19902 594
rect 19842 538 19852 578
rect 19892 538 19902 578
rect 19842 478 19902 538
rect 19842 464 19852 478
rect 19410 338 19420 378
rect 19460 338 19470 378
rect 19410 278 19470 338
rect 19410 238 19420 278
rect 19460 238 19470 278
rect 19410 32 19470 238
rect 19554 378 19614 400
rect 19554 338 19564 378
rect 19604 338 19614 378
rect 19554 278 19614 338
rect 19554 238 19564 278
rect 19604 238 19614 278
rect 19554 188 19614 238
rect 19698 378 19758 438
rect 19840 458 19852 464
rect 19892 464 19902 478
rect 19986 578 20046 594
rect 19986 538 19996 578
rect 20036 538 20046 578
rect 19986 478 20046 538
rect 19892 458 19904 464
rect 19840 406 19846 458
rect 19898 406 19904 458
rect 19840 400 19904 406
rect 19986 438 19996 478
rect 20036 438 20046 478
rect 20130 578 20190 594
rect 20130 538 20140 578
rect 20180 538 20190 578
rect 20130 478 20190 538
rect 20130 464 20140 478
rect 19698 338 19708 378
rect 19748 338 19758 378
rect 19698 278 19758 338
rect 19698 238 19708 278
rect 19748 238 19758 278
rect 19698 32 19758 238
rect 19842 378 19902 400
rect 19842 338 19852 378
rect 19892 338 19902 378
rect 19842 278 19902 338
rect 19842 238 19852 278
rect 19892 238 19902 278
rect 19842 188 19902 238
rect 19986 378 20046 438
rect 20128 458 20140 464
rect 20180 464 20190 478
rect 20274 578 20334 594
rect 20274 538 20284 578
rect 20324 538 20334 578
rect 20274 478 20334 538
rect 20180 458 20192 464
rect 20128 406 20134 458
rect 20186 406 20192 458
rect 20128 400 20192 406
rect 20274 438 20284 478
rect 20324 438 20334 478
rect 20418 578 20478 594
rect 20418 538 20428 578
rect 20468 538 20478 578
rect 20418 478 20478 538
rect 20418 464 20428 478
rect 19986 338 19996 378
rect 20036 338 20046 378
rect 19986 278 20046 338
rect 19986 238 19996 278
rect 20036 238 20046 278
rect 19986 32 20046 238
rect 20130 378 20190 400
rect 20130 338 20140 378
rect 20180 338 20190 378
rect 20130 278 20190 338
rect 20130 238 20140 278
rect 20180 238 20190 278
rect 20130 188 20190 238
rect 20274 378 20334 438
rect 20416 458 20428 464
rect 20468 464 20478 478
rect 20562 578 20622 594
rect 20562 538 20572 578
rect 20612 538 20622 578
rect 20562 478 20622 538
rect 20468 458 20480 464
rect 20416 406 20422 458
rect 20474 406 20480 458
rect 20416 400 20480 406
rect 20562 438 20572 478
rect 20612 438 20622 478
rect 20706 578 20766 594
rect 20706 538 20716 578
rect 20756 538 20766 578
rect 20706 478 20766 538
rect 20706 464 20716 478
rect 20274 338 20284 378
rect 20324 338 20334 378
rect 20274 278 20334 338
rect 20274 238 20284 278
rect 20324 238 20334 278
rect 20274 32 20334 238
rect 20418 378 20478 400
rect 20418 338 20428 378
rect 20468 338 20478 378
rect 20418 278 20478 338
rect 20418 238 20428 278
rect 20468 238 20478 278
rect 20418 188 20478 238
rect 20562 378 20622 438
rect 20704 458 20716 464
rect 20756 464 20766 478
rect 20850 578 20910 594
rect 20850 538 20860 578
rect 20900 538 20910 578
rect 20850 478 20910 538
rect 20756 458 20768 464
rect 20704 406 20710 458
rect 20762 406 20768 458
rect 20704 400 20768 406
rect 20850 438 20860 478
rect 20900 438 20910 478
rect 20562 338 20572 378
rect 20612 338 20622 378
rect 20562 278 20622 338
rect 20562 238 20572 278
rect 20612 238 20622 278
rect 20562 32 20622 238
rect 20706 378 20766 400
rect 20706 338 20716 378
rect 20756 338 20766 378
rect 20706 278 20766 338
rect 20706 238 20716 278
rect 20756 238 20766 278
rect 20706 188 20766 238
rect 20850 378 20910 438
rect 20850 338 20860 378
rect 20900 338 20910 378
rect 20850 278 20910 338
rect 20850 238 20860 278
rect 20900 238 20910 278
rect 20850 32 20910 238
rect 112 26 176 32
rect 112 -26 118 26
rect 170 -26 176 26
rect 112 -32 176 -26
rect 400 26 464 32
rect 400 -26 406 26
rect 458 -26 464 26
rect 400 -32 464 -26
rect 688 26 752 32
rect 688 -26 694 26
rect 746 -26 752 26
rect 688 -32 752 -26
rect 976 26 1040 32
rect 976 -26 982 26
rect 1034 -26 1040 26
rect 976 -32 1040 -26
rect 1264 26 1328 32
rect 1264 -26 1270 26
rect 1322 -26 1328 26
rect 1264 -32 1328 -26
rect 1552 26 1616 32
rect 1552 -26 1558 26
rect 1610 -26 1616 26
rect 1552 -32 1616 -26
rect 3568 26 3632 32
rect 3568 -26 3574 26
rect 3626 -26 3632 26
rect 3568 -32 3632 -26
rect 3856 26 3920 32
rect 3856 -26 3862 26
rect 3914 -26 3920 26
rect 3856 -32 3920 -26
rect 4144 26 4208 32
rect 4144 -26 4150 26
rect 4202 -26 4208 26
rect 4144 -32 4208 -26
rect 4432 26 4496 32
rect 4432 -26 4438 26
rect 4490 -26 4496 26
rect 4432 -32 4496 -26
rect 4720 26 4784 32
rect 4720 -26 4726 26
rect 4778 -26 4784 26
rect 4720 -32 4784 -26
rect 5008 26 5072 32
rect 5008 -26 5014 26
rect 5066 -26 5072 26
rect 5008 -32 5072 -26
rect 5296 26 5360 32
rect 5296 -26 5302 26
rect 5354 -26 5360 26
rect 5296 -32 5360 -26
rect 5584 26 5648 32
rect 5584 -26 5590 26
rect 5642 -26 5648 26
rect 5584 -32 5648 -26
rect 5872 26 5936 32
rect 5872 -26 5878 26
rect 5930 -26 5936 26
rect 5872 -32 5936 -26
rect 6160 26 6224 32
rect 6160 -26 6166 26
rect 6218 -26 6224 26
rect 6160 -32 6224 -26
rect 6448 26 6512 32
rect 6448 -26 6454 26
rect 6506 -26 6512 26
rect 6448 -32 6512 -26
rect 6736 26 6800 32
rect 6736 -26 6742 26
rect 6794 -26 6800 26
rect 6736 -32 6800 -26
rect 7024 26 7088 32
rect 7024 -26 7030 26
rect 7082 -26 7088 26
rect 7024 -32 7088 -26
rect 7312 26 7376 32
rect 7312 -26 7318 26
rect 7370 -26 7376 26
rect 7312 -32 7376 -26
rect 8176 26 8240 32
rect 8176 -26 8182 26
rect 8234 -26 8240 26
rect 8176 -32 8240 -26
rect 8752 26 8816 32
rect 8752 -26 8758 26
rect 8810 -26 8816 26
rect 8752 -32 8816 -26
rect 9040 26 9104 32
rect 9040 -26 9046 26
rect 9098 -26 9104 26
rect 9040 -32 9104 -26
rect 9328 26 9392 32
rect 9328 -26 9334 26
rect 9386 -26 9392 26
rect 9328 -32 9392 -26
rect 9616 26 9680 32
rect 9616 -26 9622 26
rect 9674 -26 9680 26
rect 9616 -32 9680 -26
rect 9904 26 9968 32
rect 9904 -26 9910 26
rect 9962 -26 9968 26
rect 9904 -32 9968 -26
rect 10192 26 10256 32
rect 10192 -26 10198 26
rect 10250 -26 10256 26
rect 10192 -32 10256 -26
rect 11056 26 11120 32
rect 11056 -26 11062 26
rect 11114 -26 11120 26
rect 11056 -32 11120 -26
rect 11920 26 11984 32
rect 11920 -26 11926 26
rect 11978 -26 11984 26
rect 11920 -32 11984 -26
rect 12208 26 12272 32
rect 12208 -26 12214 26
rect 12266 -26 12272 26
rect 12208 -32 12272 -26
rect 12496 26 12560 32
rect 12496 -26 12502 26
rect 12554 -26 12560 26
rect 12496 -32 12560 -26
rect 12784 26 12848 32
rect 12784 -26 12790 26
rect 12842 -26 12848 26
rect 12784 -32 12848 -26
rect 13072 26 13136 32
rect 13072 -26 13078 26
rect 13130 -26 13136 26
rect 13072 -32 13136 -26
rect 13360 26 13424 32
rect 13360 -26 13366 26
rect 13418 -26 13424 26
rect 13360 -32 13424 -26
rect 13648 26 13712 32
rect 13648 -26 13654 26
rect 13706 -26 13712 26
rect 13648 -32 13712 -26
rect 13936 26 14000 32
rect 13936 -26 13942 26
rect 13994 -26 14000 26
rect 13936 -32 14000 -26
rect 14224 26 14288 32
rect 14224 -26 14230 26
rect 14282 -26 14288 26
rect 14224 -32 14288 -26
rect 14512 26 14576 32
rect 14512 -26 14518 26
rect 14570 -26 14576 26
rect 14512 -32 14576 -26
rect 14800 26 14864 32
rect 14800 -26 14806 26
rect 14858 -26 14864 26
rect 14800 -32 14864 -26
rect 15088 26 15152 32
rect 15088 -26 15094 26
rect 15146 -26 15152 26
rect 15088 -32 15152 -26
rect 15376 26 15440 32
rect 15376 -26 15382 26
rect 15434 -26 15440 26
rect 15376 -32 15440 -26
rect 15664 26 15728 32
rect 15664 -26 15670 26
rect 15722 -26 15728 26
rect 15664 -32 15728 -26
rect 15952 26 16016 32
rect 15952 -26 15958 26
rect 16010 -26 16016 26
rect 15952 -32 16016 -26
rect 16240 26 16304 32
rect 16240 -26 16246 26
rect 16298 -26 16304 26
rect 16240 -32 16304 -26
rect 16528 26 16592 32
rect 16528 -26 16534 26
rect 16586 -26 16592 26
rect 16528 -32 16592 -26
rect 16816 26 16880 32
rect 16816 -26 16822 26
rect 16874 -26 16880 26
rect 16816 -32 16880 -26
rect 17104 26 17168 32
rect 17104 -26 17110 26
rect 17162 -26 17168 26
rect 17104 -32 17168 -26
rect 17392 26 17456 32
rect 17392 -26 17398 26
rect 17450 -26 17456 26
rect 17392 -32 17456 -26
rect 17680 26 17744 32
rect 17680 -26 17686 26
rect 17738 -26 17744 26
rect 17680 -32 17744 -26
rect 17968 26 18032 32
rect 17968 -26 17974 26
rect 18026 -26 18032 26
rect 17968 -32 18032 -26
rect 18256 26 18320 32
rect 18256 -26 18262 26
rect 18314 -26 18320 26
rect 18256 -32 18320 -26
rect 18544 26 18608 32
rect 18544 -26 18550 26
rect 18602 -26 18608 26
rect 18544 -32 18608 -26
rect 18832 26 18896 32
rect 18832 -26 18838 26
rect 18890 -26 18896 26
rect 18832 -32 18896 -26
rect 19120 26 19184 32
rect 19120 -26 19126 26
rect 19178 -26 19184 26
rect 19120 -32 19184 -26
rect 19408 26 19472 32
rect 19408 -26 19414 26
rect 19466 -26 19472 26
rect 19408 -32 19472 -26
rect 19696 26 19760 32
rect 19696 -26 19702 26
rect 19754 -26 19760 26
rect 19696 -32 19760 -26
rect 19984 26 20048 32
rect 19984 -26 19990 26
rect 20042 -26 20048 26
rect 19984 -32 20048 -26
rect 20272 26 20336 32
rect 20272 -26 20278 26
rect 20330 -26 20336 26
rect 20272 -32 20336 -26
rect 20560 26 20624 32
rect 20560 -26 20566 26
rect 20618 -26 20624 26
rect 20560 -32 20624 -26
rect 20848 26 20912 32
rect 20848 -26 20854 26
rect 20906 -26 20912 26
rect 20848 -32 20912 -26
rect 114 -40 174 -32
rect 402 -40 462 -32
rect 690 -40 750 -32
rect 978 -40 1038 -32
rect 1266 -40 1326 -32
rect 1554 -40 1614 -32
rect 3570 -40 3630 -32
rect 3858 -40 3918 -32
rect 4146 -40 4206 -32
rect 4434 -40 4494 -32
rect 4722 -40 4782 -32
rect 5010 -40 5070 -32
rect 5298 -40 5358 -32
rect 5586 -40 5646 -32
rect 5874 -40 5934 -32
rect 6162 -40 6222 -32
rect 6450 -40 6510 -32
rect 6738 -40 6798 -32
rect 7026 -40 7086 -32
rect 7314 -40 7374 -32
rect 8754 -40 8814 -32
rect 9042 -40 9102 -32
rect 9330 -40 9390 -32
rect 9618 -40 9678 -32
rect 9906 -40 9966 -32
rect 10194 -40 10254 -32
rect 11922 -40 11982 -32
rect 12210 -40 12270 -32
rect 12498 -40 12558 -32
rect 12786 -40 12846 -32
rect 13074 -40 13134 -32
rect 13362 -40 13422 -32
rect 13650 -40 13710 -32
rect 13938 -40 13998 -32
rect 14226 -40 14286 -32
rect 14514 -40 14574 -32
rect 14802 -40 14862 -32
rect 15090 -40 15150 -32
rect 15378 -40 15438 -32
rect 15666 -40 15726 -32
rect 15954 -40 16014 -32
rect 16242 -40 16302 -32
rect 16530 -40 16590 -32
rect 16818 -40 16878 -32
rect 17106 -40 17166 -32
rect 17394 -40 17454 -32
rect 17682 -40 17742 -32
rect 17970 -40 18030 -32
rect 18258 -40 18318 -32
rect 18546 -40 18606 -32
rect 18834 -40 18894 -32
rect 19122 -40 19182 -32
rect 19410 -40 19470 -32
rect 19698 -40 19758 -32
rect 19986 -40 20046 -32
rect 20274 -40 20334 -32
rect 20562 -40 20622 -32
rect 20850 -40 20910 -32
<< via1 >>
rect 118 4006 170 4058
rect 406 4006 458 4058
rect 694 4006 746 4058
rect 982 4006 1034 4058
rect 1270 4006 1322 4058
rect 1558 4006 1610 4058
rect 1846 4006 1898 4058
rect 2134 4006 2186 4058
rect 2422 4006 2474 4058
rect 2710 4006 2762 4058
rect 2998 4006 3050 4058
rect 3286 4006 3338 4058
rect 3574 4006 3626 4058
rect 3862 4006 3914 4058
rect 4150 4006 4202 4058
rect 4438 4006 4490 4058
rect 4726 4006 4778 4058
rect 5014 4006 5066 4058
rect 5302 4006 5354 4058
rect 5590 4006 5642 4058
rect 6454 4006 6506 4058
rect 7030 4006 7082 4058
rect 7318 4006 7370 4058
rect 7606 4006 7658 4058
rect 7894 4006 7946 4058
rect 8182 4006 8234 4058
rect 8470 4006 8522 4058
rect 9334 4006 9386 4058
rect 10198 4006 10250 4058
rect 10486 4006 10538 4058
rect 10774 4006 10826 4058
rect 11062 4006 11114 4058
rect 11350 4006 11402 4058
rect 11638 4006 11690 4058
rect 11926 4006 11978 4058
rect 12214 4006 12266 4058
rect 14230 4006 14282 4058
rect 14518 4006 14570 4058
rect 14806 4006 14858 4058
rect 15094 4006 15146 4058
rect 15382 4006 15434 4058
rect 15670 4006 15722 4058
rect 15958 4006 16010 4058
rect 16246 4006 16298 4058
rect 16534 4006 16586 4058
rect 16822 4006 16874 4058
rect 17110 4006 17162 4058
rect 17398 4006 17450 4058
rect 17686 4006 17738 4058
rect 17974 4006 18026 4058
rect 18262 4006 18314 4058
rect 18550 4006 18602 4058
rect 18838 4006 18890 4058
rect 19126 4006 19178 4058
rect 19414 4006 19466 4058
rect 19702 4006 19754 4058
rect 19990 4006 20042 4058
rect 262 3574 268 3626
rect 268 3574 308 3626
rect 308 3574 314 3626
rect 838 3594 890 3626
rect 838 3574 844 3594
rect 844 3574 884 3594
rect 884 3574 890 3594
rect 1414 3594 1466 3626
rect 1414 3574 1420 3594
rect 1420 3574 1460 3594
rect 1460 3574 1466 3594
rect 1990 3594 2042 3626
rect 1990 3574 1996 3594
rect 1996 3574 2036 3594
rect 2036 3574 2042 3594
rect 2566 3594 2618 3626
rect 2566 3574 2572 3594
rect 2572 3574 2612 3594
rect 2612 3574 2618 3594
rect 3142 3594 3194 3626
rect 3142 3574 3148 3594
rect 3148 3574 3188 3594
rect 3188 3574 3194 3594
rect 3718 3574 3724 3626
rect 3724 3574 3764 3626
rect 3764 3574 3770 3626
rect 4294 3594 4346 3626
rect 4294 3574 4300 3594
rect 4300 3574 4340 3594
rect 4340 3574 4346 3594
rect 4870 3594 4922 3626
rect 4870 3574 4876 3594
rect 4876 3574 4916 3594
rect 4916 3574 4922 3594
rect 5446 3594 5498 3626
rect 5446 3574 5452 3594
rect 5452 3574 5492 3594
rect 5492 3574 5498 3594
rect 6022 3754 6028 3770
rect 6028 3754 6068 3770
rect 6068 3754 6074 3770
rect 6022 3718 6074 3754
rect 5878 3594 5930 3626
rect 5878 3574 5884 3594
rect 5884 3574 5924 3594
rect 5924 3574 5930 3594
rect 6166 3594 6218 3626
rect 6166 3574 6172 3594
rect 6172 3574 6212 3594
rect 6212 3574 6218 3594
rect 6742 3754 6748 3770
rect 6748 3754 6788 3770
rect 6788 3754 6794 3770
rect 6742 3718 6794 3754
rect 7174 3574 7180 3626
rect 7180 3574 7220 3626
rect 7220 3574 7226 3626
rect 7750 3594 7802 3626
rect 7750 3574 7756 3594
rect 7756 3574 7796 3594
rect 7796 3574 7802 3594
rect 8326 3594 8378 3626
rect 8326 3574 8332 3594
rect 8332 3574 8372 3594
rect 8372 3574 8378 3594
rect 8902 3754 8908 3770
rect 8908 3754 8948 3770
rect 8948 3754 8954 3770
rect 8902 3718 8954 3754
rect 8758 3594 8810 3626
rect 8758 3574 8764 3594
rect 8764 3574 8804 3594
rect 8804 3574 8810 3594
rect 9046 3594 9098 3626
rect 9046 3574 9052 3594
rect 9052 3574 9092 3594
rect 9092 3574 9098 3594
rect 9622 3754 9628 3770
rect 9628 3754 9668 3770
rect 9668 3754 9674 3770
rect 9622 3718 9674 3754
rect 10342 3594 10394 3626
rect 10342 3574 10348 3594
rect 10348 3574 10388 3594
rect 10388 3574 10394 3594
rect 10918 3594 10970 3626
rect 10918 3574 10924 3594
rect 10924 3574 10964 3594
rect 10964 3574 10970 3594
rect 11494 3574 11500 3626
rect 11500 3574 11540 3626
rect 11540 3574 11546 3626
rect 12502 3754 12508 3770
rect 12508 3754 12548 3770
rect 12548 3754 12554 3770
rect 12502 3718 12554 3754
rect 12070 3594 12122 3626
rect 12070 3574 12076 3594
rect 12076 3574 12116 3594
rect 12116 3574 12122 3594
rect 12790 3754 12796 3770
rect 12796 3754 12836 3770
rect 12836 3754 12842 3770
rect 12790 3718 12842 3754
rect 13654 3754 13660 3770
rect 13660 3754 13700 3770
rect 13700 3754 13706 3770
rect 13654 3718 13706 3754
rect 12646 3594 12698 3626
rect 12646 3574 12652 3594
rect 12652 3574 12692 3594
rect 12692 3574 12698 3594
rect 13942 3754 13948 3770
rect 13948 3754 13988 3770
rect 13988 3754 13994 3770
rect 13942 3718 13994 3754
rect 13798 3594 13850 3626
rect 13798 3574 13804 3594
rect 13804 3574 13844 3594
rect 13844 3574 13850 3594
rect 14374 3594 14426 3626
rect 14374 3574 14380 3594
rect 14380 3574 14420 3594
rect 14420 3574 14426 3594
rect 14950 3594 15002 3626
rect 14950 3574 14956 3594
rect 14956 3574 14996 3594
rect 14996 3574 15002 3594
rect 15526 3574 15532 3626
rect 15532 3574 15572 3626
rect 15572 3574 15578 3626
rect 16102 3574 16108 3626
rect 16108 3574 16148 3626
rect 16148 3574 16154 3626
rect 16678 3594 16730 3626
rect 16678 3574 16684 3594
rect 16684 3574 16724 3594
rect 16724 3574 16730 3594
rect 16966 3594 17018 3626
rect 16966 3574 16972 3594
rect 16972 3574 17012 3594
rect 17012 3574 17018 3594
rect 17254 3594 17306 3626
rect 17254 3574 17260 3594
rect 17260 3574 17300 3594
rect 17300 3574 17306 3594
rect 17542 3594 17594 3626
rect 17542 3574 17548 3594
rect 17548 3574 17588 3594
rect 17588 3574 17594 3594
rect 17830 3594 17882 3626
rect 17830 3574 17836 3594
rect 17836 3574 17876 3594
rect 17876 3574 17882 3594
rect 18118 3594 18170 3626
rect 18118 3574 18124 3594
rect 18124 3574 18164 3594
rect 18164 3574 18170 3594
rect 18406 3594 18458 3626
rect 18406 3574 18412 3594
rect 18412 3574 18452 3594
rect 18452 3574 18458 3594
rect 18694 3594 18746 3626
rect 18694 3574 18700 3594
rect 18700 3574 18740 3594
rect 18740 3574 18746 3594
rect 18982 3594 19034 3626
rect 18982 3574 18988 3594
rect 18988 3574 19028 3594
rect 19028 3574 19034 3594
rect 19270 3594 19322 3626
rect 19270 3574 19276 3594
rect 19276 3574 19316 3594
rect 19316 3574 19322 3594
rect 19558 3594 19610 3626
rect 19558 3574 19564 3594
rect 19564 3574 19604 3594
rect 19604 3574 19610 3594
rect 19846 3594 19898 3626
rect 19846 3574 19852 3594
rect 19852 3574 19892 3594
rect 19892 3574 19898 3594
rect 838 3286 890 3338
rect 1414 3286 1466 3338
rect 1990 3286 2042 3338
rect 2566 3286 2618 3338
rect 3142 3286 3194 3338
rect 4294 3286 4346 3338
rect 4870 3286 4922 3338
rect 5446 3286 5498 3338
rect 6022 3286 6074 3338
rect 6742 3330 6794 3338
rect 6742 3294 6752 3330
rect 6752 3294 6788 3330
rect 6788 3294 6794 3330
rect 6742 3286 6794 3294
rect 7750 3286 7802 3338
rect 8326 3286 8378 3338
rect 8902 3286 8954 3338
rect 9622 3330 9674 3338
rect 9622 3294 9632 3330
rect 9632 3294 9668 3330
rect 9668 3294 9674 3330
rect 9622 3286 9674 3294
rect 10342 3286 10394 3338
rect 10918 3286 10970 3338
rect 12070 3286 12122 3338
rect 12646 3286 12698 3338
rect 13798 3286 13850 3338
rect 14374 3286 14426 3338
rect 14950 3286 15002 3338
rect 16678 3286 16730 3338
rect 16966 3286 17018 3338
rect 17254 3286 17306 3338
rect 17542 3286 17594 3338
rect 17830 3286 17882 3338
rect 18118 3286 18170 3338
rect 18406 3286 18458 3338
rect 18694 3286 18746 3338
rect 18982 3286 19034 3338
rect 19270 3286 19322 3338
rect 19558 3286 19610 3338
rect 19846 3286 19898 3338
rect 6454 2998 6506 3050
rect 9334 2998 9386 3050
rect 838 2710 890 2762
rect 1414 2710 1466 2762
rect 1990 2710 2042 2762
rect 2566 2710 2618 2762
rect 3142 2710 3194 2762
rect 4294 2710 4346 2762
rect 4870 2710 4922 2762
rect 5446 2710 5498 2762
rect 6022 2710 6074 2762
rect 6742 2754 6794 2762
rect 6742 2718 6746 2754
rect 6746 2718 6782 2754
rect 6782 2718 6794 2754
rect 6742 2710 6794 2718
rect 7750 2710 7802 2762
rect 8326 2710 8378 2762
rect 8902 2710 8954 2762
rect 9622 2754 9674 2762
rect 9622 2718 9626 2754
rect 9626 2718 9662 2754
rect 9662 2718 9674 2754
rect 9622 2710 9674 2718
rect 10342 2710 10394 2762
rect 10918 2710 10970 2762
rect 12070 2710 12122 2762
rect 12646 2710 12698 2762
rect 13798 2710 13850 2762
rect 14374 2710 14426 2762
rect 14950 2710 15002 2762
rect 16678 2710 16730 2762
rect 16966 2710 17018 2762
rect 17254 2710 17306 2762
rect 17542 2710 17594 2762
rect 17830 2710 17882 2762
rect 18118 2710 18170 2762
rect 18406 2710 18458 2762
rect 18694 2710 18746 2762
rect 18982 2710 19034 2762
rect 19270 2710 19322 2762
rect 19558 2710 19610 2762
rect 19846 2710 19898 2762
rect 262 2422 314 2474
rect 838 2422 890 2474
rect 1414 2422 1466 2474
rect 1990 2422 2042 2474
rect 2566 2422 2618 2474
rect 3142 2422 3194 2474
rect 3718 2422 3770 2474
rect 4294 2422 4346 2474
rect 4870 2422 4922 2474
rect 5446 2422 5498 2474
rect 5878 2422 5930 2474
rect 6166 2422 6218 2474
rect 6022 2278 6074 2330
rect 6742 2278 6794 2330
rect 7174 2422 7226 2474
rect 7750 2422 7802 2474
rect 8326 2422 8378 2474
rect 8758 2422 8810 2474
rect 9046 2422 9098 2474
rect 8902 2278 8954 2330
rect 9622 2278 9674 2330
rect 10342 2422 10394 2474
rect 10918 2422 10970 2474
rect 11494 2422 11546 2474
rect 12070 2422 12122 2474
rect 12646 2422 12698 2474
rect 12502 2278 12554 2330
rect 13798 2422 13850 2474
rect 12790 2278 12842 2330
rect 13654 2278 13706 2330
rect 13942 2278 13994 2330
rect 14374 2422 14426 2474
rect 14950 2422 15002 2474
rect 15526 2422 15578 2474
rect 16102 2422 16154 2474
rect 16678 2422 16730 2474
rect 16966 2422 17018 2474
rect 17254 2422 17306 2474
rect 17542 2422 17594 2474
rect 17830 2422 17882 2474
rect 18118 2422 18170 2474
rect 18406 2422 18458 2474
rect 18694 2422 18746 2474
rect 18982 2422 19034 2474
rect 19270 2422 19322 2474
rect 19558 2422 19610 2474
rect 19846 2422 19898 2474
rect 118 1990 170 2042
rect 406 1990 458 2042
rect 694 1990 746 2042
rect 982 1990 1034 2042
rect 1270 1990 1322 2042
rect 1558 1990 1610 2042
rect 1846 1990 1898 2042
rect 2134 1990 2186 2042
rect 2422 1990 2474 2042
rect 2710 1990 2762 2042
rect 2998 1990 3050 2042
rect 3286 1990 3338 2042
rect 3574 1990 3626 2042
rect 3862 1990 3914 2042
rect 4150 1990 4202 2042
rect 4438 1990 4490 2042
rect 4726 1990 4778 2042
rect 5014 1990 5066 2042
rect 5302 1990 5354 2042
rect 5590 1990 5642 2042
rect 5878 1990 5930 2042
rect 6166 1990 6218 2042
rect 6454 1990 6506 2042
rect 6742 1990 6794 2042
rect 7030 1990 7082 2042
rect 7318 1990 7370 2042
rect 7606 1990 7658 2042
rect 7894 1990 7946 2042
rect 8182 1990 8234 2042
rect 8470 1990 8522 2042
rect 8758 1990 8810 2042
rect 9046 1990 9098 2042
rect 9334 1990 9386 2042
rect 9622 1990 9674 2042
rect 9910 1990 9962 2042
rect 10198 1990 10250 2042
rect 10486 1990 10538 2042
rect 10774 1990 10826 2042
rect 11062 1990 11114 2042
rect 11350 1990 11402 2042
rect 11638 1990 11690 2042
rect 11926 1990 11978 2042
rect 12214 1990 12266 2042
rect 12502 1990 12554 2042
rect 12790 1990 12842 2042
rect 13078 1990 13130 2042
rect 13366 1990 13418 2042
rect 13654 1990 13706 2042
rect 13942 1990 13994 2042
rect 14230 1990 14282 2042
rect 14518 1990 14570 2042
rect 14806 1990 14858 2042
rect 15094 1990 15146 2042
rect 15382 1990 15434 2042
rect 15670 1990 15722 2042
rect 15958 1990 16010 2042
rect 16246 1990 16298 2042
rect 16534 1990 16586 2042
rect 16822 1990 16874 2042
rect 17110 1990 17162 2042
rect 17398 1990 17450 2042
rect 17686 1990 17738 2042
rect 17974 1990 18026 2042
rect 18262 1990 18314 2042
rect 18550 1990 18602 2042
rect 18838 1990 18890 2042
rect 19126 1990 19178 2042
rect 19414 1990 19466 2042
rect 19702 1990 19754 2042
rect 19990 1990 20042 2042
rect 20278 1990 20330 2042
rect 20566 1990 20618 2042
rect 20854 1990 20906 2042
rect 262 1558 314 1610
rect 838 1558 890 1610
rect 1414 1558 1466 1610
rect 1846 1702 1898 1754
rect 2134 1702 2186 1754
rect 2998 1702 3050 1754
rect 1990 1558 2042 1610
rect 3286 1702 3338 1754
rect 3142 1558 3194 1610
rect 3718 1558 3770 1610
rect 4294 1558 4346 1610
rect 4870 1558 4922 1610
rect 5446 1558 5498 1610
rect 6022 1558 6074 1610
rect 6598 1558 6650 1610
rect 7174 1558 7226 1610
rect 7750 1702 7802 1754
rect 7606 1558 7658 1610
rect 7894 1558 7946 1610
rect 8470 1702 8522 1754
rect 8902 1558 8954 1610
rect 9478 1558 9530 1610
rect 10054 1558 10106 1610
rect 10630 1702 10682 1754
rect 10486 1558 10538 1610
rect 10774 1558 10826 1610
rect 11350 1702 11402 1754
rect 12070 1558 12122 1610
rect 12646 1558 12698 1610
rect 13222 1558 13274 1610
rect 13798 1558 13850 1610
rect 14374 1558 14426 1610
rect 14950 1558 15002 1610
rect 15526 1558 15578 1610
rect 16102 1558 16154 1610
rect 16390 1558 16442 1610
rect 16966 1558 17018 1610
rect 17542 1558 17594 1610
rect 17830 1558 17882 1610
rect 18118 1558 18170 1610
rect 18406 1558 18458 1610
rect 18694 1558 18746 1610
rect 18982 1558 19034 1610
rect 19270 1558 19322 1610
rect 19558 1558 19610 1610
rect 19846 1558 19898 1610
rect 20134 1558 20186 1610
rect 20422 1558 20474 1610
rect 20710 1558 20762 1610
rect 838 1270 890 1322
rect 1414 1270 1466 1322
rect 1990 1270 2042 1322
rect 3142 1270 3194 1322
rect 3718 1270 3770 1322
rect 4294 1270 4346 1322
rect 6022 1270 6074 1322
rect 6598 1270 6650 1322
rect 7174 1270 7226 1322
rect 7750 1270 7802 1322
rect 8470 1314 8522 1322
rect 8470 1278 8474 1314
rect 8474 1278 8510 1314
rect 8510 1278 8522 1314
rect 8470 1270 8522 1278
rect 9478 1270 9530 1322
rect 10054 1270 10106 1322
rect 10630 1270 10682 1322
rect 11350 1314 11402 1322
rect 11350 1278 11354 1314
rect 11354 1278 11390 1314
rect 11390 1278 11402 1314
rect 11350 1270 11402 1278
rect 12070 1270 12122 1322
rect 12646 1270 12698 1322
rect 13222 1270 13274 1322
rect 13798 1270 13850 1322
rect 14950 1270 15002 1322
rect 15526 1270 15578 1322
rect 16102 1270 16154 1322
rect 16390 1270 16442 1322
rect 17542 1270 17594 1322
rect 17830 1270 17882 1322
rect 18118 1270 18170 1322
rect 18406 1270 18458 1322
rect 18694 1270 18746 1322
rect 18982 1270 19034 1322
rect 19270 1270 19322 1322
rect 19558 1270 19610 1322
rect 19846 1270 19898 1322
rect 20134 1270 20186 1322
rect 20422 1270 20474 1322
rect 20710 1270 20762 1322
rect 8182 982 8234 1034
rect 11062 982 11114 1034
rect 838 694 890 746
rect 1414 694 1466 746
rect 1990 694 2042 746
rect 3142 694 3194 746
rect 3718 694 3770 746
rect 4294 694 4346 746
rect 6022 694 6074 746
rect 6598 694 6650 746
rect 7174 694 7226 746
rect 7750 694 7802 746
rect 8470 738 8522 746
rect 8470 702 8480 738
rect 8480 702 8516 738
rect 8516 702 8522 738
rect 8470 694 8522 702
rect 9478 694 9530 746
rect 10054 694 10106 746
rect 10630 694 10682 746
rect 11350 738 11402 746
rect 11350 702 11360 738
rect 11360 702 11396 738
rect 11396 702 11402 738
rect 11350 694 11402 702
rect 12070 694 12122 746
rect 12646 694 12698 746
rect 13222 694 13274 746
rect 13798 694 13850 746
rect 14950 694 15002 746
rect 15526 694 15578 746
rect 16102 694 16154 746
rect 16390 694 16442 746
rect 17542 694 17594 746
rect 17830 694 17882 746
rect 18118 694 18170 746
rect 18406 694 18458 746
rect 18694 694 18746 746
rect 18982 694 19034 746
rect 19270 694 19322 746
rect 19558 694 19610 746
rect 19846 694 19898 746
rect 20134 694 20186 746
rect 20422 694 20474 746
rect 20710 694 20762 746
rect 262 406 268 458
rect 268 406 308 458
rect 308 406 314 458
rect 838 438 844 458
rect 844 438 884 458
rect 884 438 890 458
rect 838 406 890 438
rect 1414 438 1420 458
rect 1420 438 1460 458
rect 1460 438 1466 458
rect 1414 406 1466 438
rect 1990 438 1996 458
rect 1996 438 2036 458
rect 2036 438 2042 458
rect 1990 406 2042 438
rect 1846 278 1898 314
rect 1846 262 1852 278
rect 1852 262 1892 278
rect 1892 262 1898 278
rect 3142 438 3148 458
rect 3148 438 3188 458
rect 3188 438 3194 458
rect 3142 406 3194 438
rect 2134 278 2186 314
rect 2134 262 2140 278
rect 2140 262 2180 278
rect 2180 262 2186 278
rect 2998 278 3050 314
rect 2998 262 3004 278
rect 3004 262 3044 278
rect 3044 262 3050 278
rect 3718 438 3724 458
rect 3724 438 3764 458
rect 3764 438 3770 458
rect 3718 406 3770 438
rect 3286 278 3338 314
rect 3286 262 3292 278
rect 3292 262 3332 278
rect 3332 262 3338 278
rect 4294 438 4300 458
rect 4300 438 4340 458
rect 4340 438 4346 458
rect 4294 406 4346 438
rect 4870 406 4876 458
rect 4876 406 4916 458
rect 4916 406 4922 458
rect 5446 406 5452 458
rect 5452 406 5492 458
rect 5492 406 5498 458
rect 6022 438 6028 458
rect 6028 438 6068 458
rect 6068 438 6074 458
rect 6022 406 6074 438
rect 6598 438 6604 458
rect 6604 438 6644 458
rect 6644 438 6650 458
rect 6598 406 6650 438
rect 7174 438 7180 458
rect 7180 438 7220 458
rect 7220 438 7226 458
rect 7174 406 7226 438
rect 7606 438 7612 458
rect 7612 438 7652 458
rect 7652 438 7658 458
rect 7606 406 7658 438
rect 7894 438 7900 458
rect 7900 438 7940 458
rect 7940 438 7946 458
rect 7894 406 7946 438
rect 7750 278 7802 314
rect 7750 262 7756 278
rect 7756 262 7796 278
rect 7796 262 7802 278
rect 8902 406 8908 458
rect 8908 406 8948 458
rect 8948 406 8954 458
rect 8470 278 8522 314
rect 8470 262 8476 278
rect 8476 262 8516 278
rect 8516 262 8522 278
rect 9478 438 9484 458
rect 9484 438 9524 458
rect 9524 438 9530 458
rect 9478 406 9530 438
rect 10054 438 10060 458
rect 10060 438 10100 458
rect 10100 438 10106 458
rect 10054 406 10106 438
rect 10486 438 10492 458
rect 10492 438 10532 458
rect 10532 438 10538 458
rect 10486 406 10538 438
rect 10774 438 10780 458
rect 10780 438 10820 458
rect 10820 438 10826 458
rect 10774 406 10826 438
rect 10630 278 10682 314
rect 10630 262 10636 278
rect 10636 262 10676 278
rect 10676 262 10682 278
rect 12070 438 12076 458
rect 12076 438 12116 458
rect 12116 438 12122 458
rect 12070 406 12122 438
rect 11350 278 11402 314
rect 11350 262 11356 278
rect 11356 262 11396 278
rect 11396 262 11402 278
rect 12646 438 12652 458
rect 12652 438 12692 458
rect 12692 438 12698 458
rect 12646 406 12698 438
rect 13222 438 13228 458
rect 13228 438 13268 458
rect 13268 438 13274 458
rect 13222 406 13274 438
rect 13798 438 13804 458
rect 13804 438 13844 458
rect 13844 438 13850 458
rect 13798 406 13850 438
rect 14374 406 14380 458
rect 14380 406 14420 458
rect 14420 406 14426 458
rect 14950 438 14956 458
rect 14956 438 14996 458
rect 14996 438 15002 458
rect 14950 406 15002 438
rect 15526 438 15532 458
rect 15532 438 15572 458
rect 15572 438 15578 458
rect 15526 406 15578 438
rect 16102 438 16108 458
rect 16108 438 16148 458
rect 16148 438 16154 458
rect 16102 406 16154 438
rect 16390 438 16396 458
rect 16396 438 16436 458
rect 16436 438 16442 458
rect 16390 406 16442 438
rect 16966 406 16972 458
rect 16972 406 17012 458
rect 17012 406 17018 458
rect 17542 438 17548 458
rect 17548 438 17588 458
rect 17588 438 17594 458
rect 17542 406 17594 438
rect 17830 438 17836 458
rect 17836 438 17876 458
rect 17876 438 17882 458
rect 17830 406 17882 438
rect 18118 438 18124 458
rect 18124 438 18164 458
rect 18164 438 18170 458
rect 18118 406 18170 438
rect 18406 438 18412 458
rect 18412 438 18452 458
rect 18452 438 18458 458
rect 18406 406 18458 438
rect 18694 438 18700 458
rect 18700 438 18740 458
rect 18740 438 18746 458
rect 18694 406 18746 438
rect 18982 438 18988 458
rect 18988 438 19028 458
rect 19028 438 19034 458
rect 18982 406 19034 438
rect 19270 438 19276 458
rect 19276 438 19316 458
rect 19316 438 19322 458
rect 19270 406 19322 438
rect 19558 438 19564 458
rect 19564 438 19604 458
rect 19604 438 19610 458
rect 19558 406 19610 438
rect 19846 438 19852 458
rect 19852 438 19892 458
rect 19892 438 19898 458
rect 19846 406 19898 438
rect 20134 438 20140 458
rect 20140 438 20180 458
rect 20180 438 20186 458
rect 20134 406 20186 438
rect 20422 438 20428 458
rect 20428 438 20468 458
rect 20468 438 20474 458
rect 20422 406 20474 438
rect 20710 438 20716 458
rect 20716 438 20756 458
rect 20756 438 20762 458
rect 20710 406 20762 438
rect 118 -26 170 26
rect 406 -26 458 26
rect 694 -26 746 26
rect 982 -26 1034 26
rect 1270 -26 1322 26
rect 1558 -26 1610 26
rect 3574 -26 3626 26
rect 3862 -26 3914 26
rect 4150 -26 4202 26
rect 4438 -26 4490 26
rect 4726 -26 4778 26
rect 5014 -26 5066 26
rect 5302 -26 5354 26
rect 5590 -26 5642 26
rect 5878 -26 5930 26
rect 6166 -26 6218 26
rect 6454 -26 6506 26
rect 6742 -26 6794 26
rect 7030 -26 7082 26
rect 7318 -26 7370 26
rect 8182 -26 8234 26
rect 8758 -26 8810 26
rect 9046 -26 9098 26
rect 9334 -26 9386 26
rect 9622 -26 9674 26
rect 9910 -26 9962 26
rect 10198 -26 10250 26
rect 11062 -26 11114 26
rect 11926 -26 11978 26
rect 12214 -26 12266 26
rect 12502 -26 12554 26
rect 12790 -26 12842 26
rect 13078 -26 13130 26
rect 13366 -26 13418 26
rect 13654 -26 13706 26
rect 13942 -26 13994 26
rect 14230 -26 14282 26
rect 14518 -26 14570 26
rect 14806 -26 14858 26
rect 15094 -26 15146 26
rect 15382 -26 15434 26
rect 15670 -26 15722 26
rect 15958 -26 16010 26
rect 16246 -26 16298 26
rect 16534 -26 16586 26
rect 16822 -26 16874 26
rect 17110 -26 17162 26
rect 17398 -26 17450 26
rect 17686 -26 17738 26
rect 17974 -26 18026 26
rect 18262 -26 18314 26
rect 18550 -26 18602 26
rect 18838 -26 18890 26
rect 19126 -26 19178 26
rect 19414 -26 19466 26
rect 19702 -26 19754 26
rect 19990 -26 20042 26
rect 20278 -26 20330 26
rect 20566 -26 20618 26
rect 20854 -26 20906 26
<< metal2 >>
rect -40 4058 21064 4092
rect -40 4006 118 4058
rect 170 4006 406 4058
rect 458 4006 694 4058
rect 746 4006 982 4058
rect 1034 4006 1270 4058
rect 1322 4006 1558 4058
rect 1610 4006 1846 4058
rect 1898 4006 2134 4058
rect 2186 4006 2422 4058
rect 2474 4006 2710 4058
rect 2762 4006 2998 4058
rect 3050 4006 3286 4058
rect 3338 4006 3574 4058
rect 3626 4006 3862 4058
rect 3914 4006 4150 4058
rect 4202 4006 4438 4058
rect 4490 4006 4726 4058
rect 4778 4006 5014 4058
rect 5066 4006 5302 4058
rect 5354 4006 5590 4058
rect 5642 4006 6454 4058
rect 6506 4006 7030 4058
rect 7082 4006 7318 4058
rect 7370 4006 7606 4058
rect 7658 4006 7894 4058
rect 7946 4006 8182 4058
rect 8234 4006 8470 4058
rect 8522 4006 9334 4058
rect 9386 4006 10198 4058
rect 10250 4006 10486 4058
rect 10538 4006 10774 4058
rect 10826 4006 11062 4058
rect 11114 4006 11350 4058
rect 11402 4006 11638 4058
rect 11690 4006 11926 4058
rect 11978 4006 12214 4058
rect 12266 4006 14230 4058
rect 14282 4006 14518 4058
rect 14570 4006 14806 4058
rect 14858 4006 15094 4058
rect 15146 4006 15382 4058
rect 15434 4006 15670 4058
rect 15722 4006 15958 4058
rect 16010 4006 16246 4058
rect 16298 4006 16534 4058
rect 16586 4006 16822 4058
rect 16874 4006 17110 4058
rect 17162 4006 17398 4058
rect 17450 4006 17686 4058
rect 17738 4006 17974 4058
rect 18026 4006 18262 4058
rect 18314 4006 18550 4058
rect 18602 4006 18838 4058
rect 18890 4006 19126 4058
rect 19178 4006 19414 4058
rect 19466 4006 19702 4058
rect 19754 4006 19990 4058
rect 20042 4006 21064 4058
rect -40 3972 21064 4006
rect 6010 3774 6086 3782
rect 5868 3772 6228 3774
rect 5868 3716 6020 3772
rect 6076 3716 6228 3772
rect 5868 3714 6228 3716
rect 6730 3772 6806 3782
rect 8890 3774 8966 3782
rect 6730 3716 6740 3772
rect 6796 3716 6806 3772
rect 6010 3706 6086 3714
rect 6730 3706 6806 3716
rect 8748 3772 9108 3774
rect 8748 3716 8900 3772
rect 8956 3716 9108 3772
rect 8748 3714 9108 3716
rect 9610 3772 9686 3782
rect 12496 3774 12560 3776
rect 12784 3774 12848 3776
rect 13648 3774 13712 3776
rect 13930 3774 14006 3782
rect 14650 3774 14726 3782
rect 9610 3716 9620 3772
rect 9676 3716 9686 3772
rect 8890 3706 8966 3714
rect 9610 3706 9686 3716
rect 12452 3772 14726 3774
rect 12452 3770 13940 3772
rect 12452 3718 12502 3770
rect 12554 3718 12790 3770
rect 12842 3718 13654 3770
rect 13706 3718 13940 3770
rect 12452 3716 13940 3718
rect 13996 3716 14660 3772
rect 14716 3716 14726 3772
rect 12452 3714 14726 3716
rect 12496 3712 12560 3714
rect 12784 3712 12848 3714
rect 13648 3712 13712 3714
rect 13930 3706 14006 3714
rect 14650 3706 14726 3714
rect 256 3630 320 3632
rect 826 3630 902 3638
rect 1402 3630 1478 3638
rect 1978 3630 2054 3638
rect 2554 3630 2630 3638
rect 3130 3630 3206 3638
rect 3712 3630 3776 3632
rect 4282 3630 4358 3638
rect 4858 3630 4934 3638
rect 5440 3630 5504 3632
rect 5872 3630 5936 3632
rect 6160 3630 6224 3632
rect 7168 3630 7232 3632
rect 7738 3630 7814 3638
rect 8320 3630 8384 3632
rect 8752 3630 8816 3632
rect 9040 3630 9104 3632
rect 10330 3630 10406 3638
rect 10906 3630 10982 3638
rect 11488 3630 11552 3632
rect 12064 3630 12128 3632
rect 12640 3630 12704 3632
rect 12922 3630 12998 3638
rect 13498 3630 13574 3638
rect 13792 3630 13856 3632
rect 14368 3630 14432 3632
rect 14938 3630 15014 3638
rect 15520 3630 15584 3632
rect 16096 3630 16160 3632
rect 16666 3630 16742 3638
rect 16960 3630 17024 3632
rect 17248 3630 17312 3632
rect 17536 3630 17600 3632
rect 17824 3630 17888 3632
rect 18112 3630 18176 3632
rect 18400 3630 18464 3632
rect 18688 3630 18752 3632
rect 18976 3630 19040 3632
rect 19264 3630 19328 3632
rect 19552 3630 19616 3632
rect 19840 3630 19904 3632
rect 144 3626 432 3630
rect 144 3574 262 3626
rect 314 3574 432 3626
rect 144 3570 432 3574
rect 684 3628 1044 3630
rect 684 3572 836 3628
rect 892 3572 1044 3628
rect 684 3570 1044 3572
rect 1260 3628 1620 3630
rect 1260 3572 1412 3628
rect 1468 3572 1620 3628
rect 1260 3570 1620 3572
rect 1836 3628 2196 3630
rect 1836 3572 1988 3628
rect 2044 3572 2196 3628
rect 1836 3570 2196 3572
rect 2412 3628 2772 3630
rect 2412 3572 2564 3628
rect 2620 3572 2772 3628
rect 2412 3570 2772 3572
rect 2988 3628 3348 3630
rect 2988 3572 3140 3628
rect 3196 3572 3348 3628
rect 2988 3570 3348 3572
rect 3600 3626 3888 3630
rect 3600 3574 3718 3626
rect 3770 3574 3888 3626
rect 3600 3570 3888 3574
rect 4140 3628 4500 3630
rect 4140 3572 4292 3628
rect 4348 3572 4500 3628
rect 4140 3570 4500 3572
rect 4716 3628 5076 3630
rect 4716 3572 4868 3628
rect 4924 3572 5076 3628
rect 4716 3570 5076 3572
rect 5292 3626 6268 3630
rect 5292 3574 5446 3626
rect 5498 3574 5878 3626
rect 5930 3574 6166 3626
rect 6218 3574 6268 3626
rect 5292 3570 6268 3574
rect 7056 3626 7344 3630
rect 7056 3574 7174 3626
rect 7226 3574 7344 3626
rect 7056 3570 7344 3574
rect 7596 3628 7956 3630
rect 7596 3572 7748 3628
rect 7804 3572 7956 3628
rect 7596 3570 7956 3572
rect 8172 3626 9148 3630
rect 8172 3574 8326 3626
rect 8378 3574 8758 3626
rect 8810 3574 9046 3626
rect 9098 3574 9148 3626
rect 8172 3570 9148 3574
rect 10188 3628 10548 3630
rect 10188 3572 10340 3628
rect 10396 3572 10548 3628
rect 10188 3570 10548 3572
rect 10764 3628 11124 3630
rect 10764 3572 10916 3628
rect 10972 3572 11124 3628
rect 10764 3570 11124 3572
rect 11376 3626 11664 3630
rect 11376 3574 11494 3626
rect 11546 3574 11664 3626
rect 11376 3570 11664 3574
rect 11916 3626 12852 3630
rect 11916 3574 12070 3626
rect 12122 3574 12646 3626
rect 12698 3574 12852 3626
rect 11916 3570 12852 3574
rect 12922 3628 13574 3630
rect 12922 3572 12932 3628
rect 12988 3572 13508 3628
rect 13564 3572 13574 3628
rect 12922 3570 13574 3572
rect 13644 3626 14580 3630
rect 13644 3574 13798 3626
rect 13850 3574 14374 3626
rect 14426 3574 14580 3626
rect 13644 3570 14580 3574
rect 14796 3628 15156 3630
rect 14796 3572 14948 3628
rect 15004 3572 15156 3628
rect 14796 3570 15156 3572
rect 15408 3626 15696 3630
rect 15408 3574 15526 3626
rect 15578 3574 15696 3626
rect 15408 3570 15696 3574
rect 15984 3626 16272 3630
rect 15984 3574 16102 3626
rect 16154 3574 16272 3626
rect 15984 3570 16272 3574
rect 16628 3628 19948 3630
rect 16628 3572 16676 3628
rect 16732 3626 19948 3628
rect 16732 3574 16966 3626
rect 17018 3574 17254 3626
rect 17306 3574 17542 3626
rect 17594 3574 17830 3626
rect 17882 3574 18118 3626
rect 18170 3574 18406 3626
rect 18458 3574 18694 3626
rect 18746 3574 18982 3626
rect 19034 3574 19270 3626
rect 19322 3574 19558 3626
rect 19610 3574 19846 3626
rect 19898 3574 19948 3626
rect 16732 3572 19948 3574
rect 16628 3570 19948 3572
rect 256 3568 320 3570
rect 826 3562 902 3570
rect 1402 3562 1478 3570
rect 1978 3562 2054 3570
rect 2554 3562 2630 3570
rect 3130 3562 3206 3570
rect 3712 3568 3776 3570
rect 4282 3562 4358 3570
rect 4858 3562 4934 3570
rect 5440 3568 5504 3570
rect 5872 3568 5936 3570
rect 6160 3568 6224 3570
rect 7168 3568 7232 3570
rect 7738 3562 7814 3570
rect 8320 3568 8384 3570
rect 8752 3568 8816 3570
rect 9040 3568 9104 3570
rect 10330 3562 10406 3570
rect 10906 3562 10982 3570
rect 11488 3568 11552 3570
rect 12064 3568 12128 3570
rect 12640 3568 12704 3570
rect 12922 3562 12998 3570
rect 13498 3562 13574 3570
rect 13792 3568 13856 3570
rect 14368 3568 14432 3570
rect 14938 3562 15014 3570
rect 15520 3568 15584 3570
rect 16096 3568 16160 3570
rect 16666 3562 16742 3570
rect 16960 3568 17024 3570
rect 17248 3568 17312 3570
rect 17536 3568 17600 3570
rect 17824 3568 17888 3570
rect 18112 3568 18176 3570
rect 18400 3568 18464 3570
rect 18688 3568 18752 3570
rect 18976 3568 19040 3570
rect 19264 3568 19328 3570
rect 19552 3568 19616 3570
rect 19840 3568 19904 3570
rect 832 3342 896 3344
rect 970 3342 1046 3350
rect 1408 3342 1472 3344
rect 1546 3342 1622 3350
rect 1984 3342 2048 3344
rect 2122 3342 2198 3350
rect 2560 3342 2624 3344
rect 2698 3342 2774 3350
rect 684 3340 1046 3342
rect 684 3338 980 3340
rect 684 3286 838 3338
rect 890 3286 980 3338
rect 684 3284 980 3286
rect 1036 3284 1046 3340
rect 684 3282 1046 3284
rect 1260 3340 1622 3342
rect 1260 3338 1556 3340
rect 1260 3286 1414 3338
rect 1466 3286 1556 3338
rect 1260 3284 1556 3286
rect 1612 3284 1622 3340
rect 1260 3282 1622 3284
rect 1836 3340 2198 3342
rect 1836 3338 2132 3340
rect 1836 3286 1990 3338
rect 2042 3286 2132 3338
rect 1836 3284 2132 3286
rect 2188 3284 2198 3340
rect 1836 3282 2198 3284
rect 2412 3340 2774 3342
rect 2412 3338 2708 3340
rect 2412 3286 2566 3338
rect 2618 3286 2708 3338
rect 2412 3284 2708 3286
rect 2764 3284 2774 3340
rect 2412 3282 2774 3284
rect 832 3280 896 3282
rect 970 3274 1046 3282
rect 1408 3280 1472 3282
rect 1546 3274 1622 3282
rect 1984 3280 2048 3282
rect 2122 3274 2198 3282
rect 2560 3280 2624 3282
rect 2698 3274 2774 3282
rect 2986 3342 3062 3350
rect 3136 3342 3200 3344
rect 4138 3342 4214 3350
rect 4288 3342 4352 3344
rect 4714 3342 4790 3350
rect 4864 3342 4928 3344
rect 5434 3342 5510 3350
rect 5866 3342 5942 3350
rect 6016 3342 6080 3344
rect 6586 3342 6662 3350
rect 6736 3342 6800 3344
rect 2986 3340 3348 3342
rect 2986 3284 2996 3340
rect 3052 3338 3348 3340
rect 3052 3286 3142 3338
rect 3194 3286 3348 3338
rect 3052 3284 3348 3286
rect 2986 3282 3348 3284
rect 4138 3340 4500 3342
rect 4138 3284 4148 3340
rect 4204 3338 4500 3340
rect 4204 3286 4294 3338
rect 4346 3286 4500 3338
rect 4204 3284 4500 3286
rect 4138 3282 4500 3284
rect 4714 3340 5076 3342
rect 4714 3284 4724 3340
rect 4780 3338 5076 3340
rect 4780 3286 4870 3338
rect 4922 3286 5076 3338
rect 4780 3284 5076 3286
rect 4714 3282 5076 3284
rect 5292 3340 5652 3342
rect 5292 3284 5444 3340
rect 5500 3284 5652 3340
rect 5292 3282 5652 3284
rect 5866 3340 6228 3342
rect 5866 3284 5876 3340
rect 5932 3338 6228 3340
rect 5932 3286 6022 3338
rect 6074 3286 6228 3338
rect 5932 3284 6228 3286
rect 5866 3282 6228 3284
rect 6586 3340 6800 3342
rect 6586 3284 6596 3340
rect 6652 3338 6800 3340
rect 6652 3286 6742 3338
rect 6794 3286 6800 3338
rect 6652 3284 6800 3286
rect 6586 3282 6800 3284
rect 2986 3274 3062 3282
rect 3136 3280 3200 3282
rect 4138 3274 4214 3282
rect 4288 3280 4352 3282
rect 4714 3274 4790 3282
rect 4864 3280 4928 3282
rect 5434 3274 5510 3282
rect 5866 3274 5942 3282
rect 6016 3280 6080 3282
rect 6586 3274 6662 3282
rect 6736 3280 6800 3282
rect 7594 3342 7670 3350
rect 7744 3342 7808 3344
rect 8314 3342 8390 3350
rect 8746 3342 8822 3350
rect 8896 3342 8960 3344
rect 9466 3342 9542 3350
rect 9616 3342 9680 3344
rect 7594 3340 7956 3342
rect 7594 3284 7604 3340
rect 7660 3338 7956 3340
rect 7660 3286 7750 3338
rect 7802 3286 7956 3338
rect 7660 3284 7956 3286
rect 7594 3282 7956 3284
rect 8172 3340 8532 3342
rect 8172 3284 8324 3340
rect 8380 3284 8532 3340
rect 8172 3282 8532 3284
rect 8746 3340 9108 3342
rect 8746 3284 8756 3340
rect 8812 3338 9108 3340
rect 8812 3286 8902 3338
rect 8954 3286 9108 3338
rect 8812 3284 9108 3286
rect 8746 3282 9108 3284
rect 9466 3340 9680 3342
rect 9466 3284 9476 3340
rect 9532 3338 9680 3340
rect 9532 3286 9622 3338
rect 9674 3286 9680 3338
rect 9532 3284 9680 3286
rect 9466 3282 9680 3284
rect 7594 3274 7670 3282
rect 7744 3280 7808 3282
rect 8314 3274 8390 3282
rect 8746 3274 8822 3282
rect 8896 3280 8960 3282
rect 9466 3274 9542 3282
rect 9616 3280 9680 3282
rect 10186 3342 10262 3350
rect 10336 3342 10400 3344
rect 10762 3342 10838 3350
rect 10912 3342 10976 3344
rect 12058 3342 12134 3350
rect 12640 3342 12704 3344
rect 12922 3342 12998 3350
rect 10186 3340 10548 3342
rect 10186 3284 10196 3340
rect 10252 3338 10548 3340
rect 10252 3286 10342 3338
rect 10394 3286 10548 3338
rect 10252 3284 10548 3286
rect 10186 3282 10548 3284
rect 10762 3340 11124 3342
rect 10762 3284 10772 3340
rect 10828 3338 11124 3340
rect 10828 3286 10918 3338
rect 10970 3286 11124 3338
rect 10828 3284 11124 3286
rect 10762 3282 11124 3284
rect 11916 3340 12276 3342
rect 11916 3284 12068 3340
rect 12124 3284 12276 3340
rect 11916 3282 12276 3284
rect 12492 3340 12998 3342
rect 12492 3338 12932 3340
rect 12492 3286 12646 3338
rect 12698 3286 12932 3338
rect 12492 3284 12932 3286
rect 12988 3284 12998 3340
rect 12492 3282 12998 3284
rect 10186 3274 10262 3282
rect 10336 3280 10400 3282
rect 10762 3274 10838 3282
rect 10912 3280 10976 3282
rect 12058 3274 12134 3282
rect 12640 3280 12704 3282
rect 12922 3274 12998 3282
rect 13210 3342 13286 3350
rect 13792 3342 13856 3344
rect 14362 3342 14438 3350
rect 14650 3342 14726 3350
rect 14944 3342 15008 3344
rect 16672 3342 16736 3344
rect 16960 3342 17024 3344
rect 17248 3342 17312 3344
rect 17536 3342 17600 3344
rect 17824 3342 17888 3344
rect 18112 3342 18176 3344
rect 18400 3342 18464 3344
rect 18688 3342 18752 3344
rect 18976 3342 19040 3344
rect 19264 3342 19328 3344
rect 19552 3342 19616 3344
rect 19840 3342 19904 3344
rect 19978 3342 20054 3350
rect 13210 3340 14004 3342
rect 13210 3284 13220 3340
rect 13276 3338 14004 3340
rect 13276 3286 13798 3338
rect 13850 3286 14004 3338
rect 13276 3284 14004 3286
rect 13210 3282 14004 3284
rect 14220 3340 14580 3342
rect 14220 3284 14372 3340
rect 14428 3284 14580 3340
rect 14220 3282 14580 3284
rect 14650 3340 15156 3342
rect 14650 3284 14660 3340
rect 14716 3338 15156 3340
rect 14716 3286 14950 3338
rect 15002 3286 15156 3338
rect 14716 3284 15156 3286
rect 14650 3282 15156 3284
rect 16628 3340 20054 3342
rect 16628 3338 19988 3340
rect 16628 3286 16678 3338
rect 16730 3286 16966 3338
rect 17018 3286 17254 3338
rect 17306 3286 17542 3338
rect 17594 3286 17830 3338
rect 17882 3286 18118 3338
rect 18170 3286 18406 3338
rect 18458 3286 18694 3338
rect 18746 3286 18982 3338
rect 19034 3286 19270 3338
rect 19322 3286 19558 3338
rect 19610 3286 19846 3338
rect 19898 3286 19988 3338
rect 16628 3284 19988 3286
rect 20044 3284 20054 3340
rect 16628 3282 20054 3284
rect 13210 3274 13286 3282
rect 13792 3280 13856 3282
rect 14362 3274 14438 3282
rect 14650 3274 14726 3282
rect 14944 3280 15008 3282
rect 16672 3280 16736 3282
rect 16960 3280 17024 3282
rect 17248 3280 17312 3282
rect 17536 3280 17600 3282
rect 17824 3280 17888 3282
rect 18112 3280 18176 3282
rect 18400 3280 18464 3282
rect 18688 3280 18752 3282
rect 18976 3280 19040 3282
rect 19264 3280 19328 3282
rect 19552 3280 19616 3282
rect 19840 3280 19904 3282
rect 19978 3274 20054 3282
rect 1546 3054 1622 3062
rect 1978 3054 2054 3062
rect 1546 3052 2054 3054
rect 1546 2996 1556 3052
rect 1612 2996 1988 3052
rect 2044 2996 2054 3052
rect 1546 2994 2054 2996
rect 1546 2986 1622 2994
rect 1978 2986 2054 2994
rect 6442 3054 6518 3062
rect 7738 3054 7814 3062
rect 8314 3054 8390 3062
rect 6442 3052 8390 3054
rect 6442 2996 6452 3052
rect 6508 2996 7748 3052
rect 7804 2996 8324 3052
rect 8380 2996 8390 3052
rect 6442 2994 8390 2996
rect 6442 2986 6518 2994
rect 7738 2986 7814 2994
rect 8314 2986 8390 2994
rect 9322 3054 9398 3062
rect 9322 3052 9668 3054
rect 9322 2996 9332 3052
rect 9388 2996 9668 3052
rect 9322 2994 9668 2996
rect 9322 2986 9398 2994
rect 832 2766 896 2768
rect 970 2766 1046 2774
rect 1408 2766 1472 2768
rect 1546 2766 1622 2774
rect 1984 2766 2048 2768
rect 2122 2766 2198 2774
rect 2560 2766 2624 2768
rect 2698 2766 2774 2774
rect 684 2764 1046 2766
rect 684 2762 980 2764
rect 684 2710 838 2762
rect 890 2710 980 2762
rect 684 2708 980 2710
rect 1036 2708 1046 2764
rect 684 2706 1046 2708
rect 1260 2764 1622 2766
rect 1260 2762 1556 2764
rect 1260 2710 1414 2762
rect 1466 2710 1556 2762
rect 1260 2708 1556 2710
rect 1612 2708 1622 2764
rect 1260 2706 1622 2708
rect 1836 2764 2198 2766
rect 1836 2762 2132 2764
rect 1836 2710 1990 2762
rect 2042 2710 2132 2762
rect 1836 2708 2132 2710
rect 2188 2708 2198 2764
rect 1836 2706 2198 2708
rect 2412 2764 2774 2766
rect 2412 2762 2708 2764
rect 2412 2710 2566 2762
rect 2618 2710 2708 2762
rect 2412 2708 2708 2710
rect 2764 2708 2774 2764
rect 2412 2706 2774 2708
rect 832 2704 896 2706
rect 970 2698 1046 2706
rect 1408 2704 1472 2706
rect 1546 2698 1622 2706
rect 1984 2704 2048 2706
rect 2122 2698 2198 2706
rect 2560 2704 2624 2706
rect 2698 2698 2774 2706
rect 2986 2766 3062 2774
rect 3136 2766 3200 2768
rect 4138 2766 4214 2774
rect 4288 2766 4352 2768
rect 4714 2766 4790 2774
rect 4864 2766 4928 2768
rect 5434 2766 5510 2774
rect 6016 2766 6080 2768
rect 6154 2766 6230 2774
rect 2986 2764 3348 2766
rect 2986 2708 2996 2764
rect 3052 2762 3348 2764
rect 3052 2710 3142 2762
rect 3194 2710 3348 2762
rect 3052 2708 3348 2710
rect 2986 2706 3348 2708
rect 4138 2764 4500 2766
rect 4138 2708 4148 2764
rect 4204 2762 4500 2764
rect 4204 2710 4294 2762
rect 4346 2710 4500 2762
rect 4204 2708 4500 2710
rect 4138 2706 4500 2708
rect 4714 2764 5076 2766
rect 4714 2708 4724 2764
rect 4780 2762 5076 2764
rect 4780 2710 4870 2762
rect 4922 2710 5076 2762
rect 4780 2708 5076 2710
rect 4714 2706 5076 2708
rect 5292 2764 5652 2766
rect 5292 2708 5444 2764
rect 5500 2708 5652 2764
rect 5292 2706 5652 2708
rect 5868 2764 6230 2766
rect 5868 2762 6164 2764
rect 5868 2710 6022 2762
rect 6074 2710 6164 2762
rect 5868 2708 6164 2710
rect 6220 2708 6230 2764
rect 5868 2706 6230 2708
rect 2986 2698 3062 2706
rect 3136 2704 3200 2706
rect 4138 2698 4214 2706
rect 4288 2704 4352 2706
rect 4714 2698 4790 2706
rect 4864 2704 4928 2706
rect 5434 2698 5510 2706
rect 6016 2704 6080 2706
rect 6154 2698 6230 2706
rect 6736 2766 6800 2768
rect 6874 2766 6950 2774
rect 6736 2764 6950 2766
rect 6736 2762 6884 2764
rect 6736 2710 6742 2762
rect 6794 2710 6884 2762
rect 6736 2708 6884 2710
rect 6940 2708 6950 2764
rect 6736 2706 6950 2708
rect 6736 2704 6800 2706
rect 6874 2698 6950 2706
rect 7594 2766 7670 2774
rect 7744 2766 7808 2768
rect 8314 2766 8390 2774
rect 8896 2766 8960 2768
rect 9034 2766 9110 2774
rect 7594 2764 7956 2766
rect 7594 2708 7604 2764
rect 7660 2762 7956 2764
rect 7660 2710 7750 2762
rect 7802 2710 7956 2762
rect 7660 2708 7956 2710
rect 7594 2706 7956 2708
rect 8172 2764 8532 2766
rect 8172 2708 8324 2764
rect 8380 2708 8532 2764
rect 8172 2706 8532 2708
rect 8748 2764 9110 2766
rect 8748 2762 9044 2764
rect 8748 2710 8902 2762
rect 8954 2710 9044 2762
rect 8748 2708 9044 2710
rect 9100 2708 9110 2764
rect 8748 2706 9110 2708
rect 7594 2698 7670 2706
rect 7744 2704 7808 2706
rect 8314 2698 8390 2706
rect 8896 2704 8960 2706
rect 9034 2698 9110 2706
rect 9616 2766 9680 2768
rect 9754 2766 9830 2774
rect 9616 2764 9830 2766
rect 9616 2762 9764 2764
rect 9616 2710 9622 2762
rect 9674 2710 9764 2762
rect 9616 2708 9764 2710
rect 9820 2708 9830 2764
rect 9616 2706 9830 2708
rect 9616 2704 9680 2706
rect 9754 2698 9830 2706
rect 10186 2766 10262 2774
rect 10336 2766 10400 2768
rect 10762 2766 10838 2774
rect 10912 2766 10976 2768
rect 12058 2766 12134 2774
rect 12640 2766 12704 2768
rect 13210 2766 13286 2774
rect 10186 2764 10548 2766
rect 10186 2708 10196 2764
rect 10252 2762 10548 2764
rect 10252 2710 10342 2762
rect 10394 2710 10548 2762
rect 10252 2708 10548 2710
rect 10186 2706 10548 2708
rect 10762 2764 11124 2766
rect 10762 2708 10772 2764
rect 10828 2762 11124 2764
rect 10828 2710 10918 2762
rect 10970 2710 11124 2762
rect 10828 2708 11124 2710
rect 10762 2706 11124 2708
rect 11916 2764 12276 2766
rect 11916 2708 12068 2764
rect 12124 2708 12276 2764
rect 11916 2706 12276 2708
rect 12492 2764 13286 2766
rect 12492 2762 13220 2764
rect 12492 2710 12646 2762
rect 12698 2710 13220 2762
rect 12492 2708 13220 2710
rect 13276 2708 13286 2764
rect 12492 2706 13286 2708
rect 10186 2698 10262 2706
rect 10336 2704 10400 2706
rect 10762 2698 10838 2706
rect 10912 2704 10976 2706
rect 12058 2698 12134 2706
rect 12640 2704 12704 2706
rect 13210 2698 13286 2706
rect 13498 2766 13574 2774
rect 13792 2766 13856 2768
rect 14362 2766 14438 2774
rect 14650 2766 14726 2774
rect 14944 2766 15008 2768
rect 16672 2766 16736 2768
rect 16960 2766 17024 2768
rect 17248 2766 17312 2768
rect 17536 2766 17600 2768
rect 17824 2766 17888 2768
rect 18112 2766 18176 2768
rect 18400 2766 18464 2768
rect 18688 2766 18752 2768
rect 18976 2766 19040 2768
rect 19264 2766 19328 2768
rect 19552 2766 19616 2768
rect 19840 2766 19904 2768
rect 19978 2766 20054 2774
rect 13498 2764 14004 2766
rect 13498 2708 13508 2764
rect 13564 2762 14004 2764
rect 13564 2710 13798 2762
rect 13850 2710 14004 2762
rect 13564 2708 14004 2710
rect 13498 2706 14004 2708
rect 14220 2764 14580 2766
rect 14220 2708 14372 2764
rect 14428 2708 14580 2764
rect 14220 2706 14580 2708
rect 14650 2764 15156 2766
rect 14650 2708 14660 2764
rect 14716 2762 15156 2764
rect 14716 2710 14950 2762
rect 15002 2710 15156 2762
rect 14716 2708 15156 2710
rect 14650 2706 15156 2708
rect 16628 2764 20054 2766
rect 16628 2762 19988 2764
rect 16628 2710 16678 2762
rect 16730 2710 16966 2762
rect 17018 2710 17254 2762
rect 17306 2710 17542 2762
rect 17594 2710 17830 2762
rect 17882 2710 18118 2762
rect 18170 2710 18406 2762
rect 18458 2710 18694 2762
rect 18746 2710 18982 2762
rect 19034 2710 19270 2762
rect 19322 2710 19558 2762
rect 19610 2710 19846 2762
rect 19898 2710 19988 2762
rect 16628 2708 19988 2710
rect 20044 2708 20054 2764
rect 16628 2706 20054 2708
rect 13498 2698 13574 2706
rect 13792 2704 13856 2706
rect 14362 2698 14438 2706
rect 14650 2698 14726 2706
rect 14944 2704 15008 2706
rect 16672 2704 16736 2706
rect 16960 2704 17024 2706
rect 17248 2704 17312 2706
rect 17536 2704 17600 2706
rect 17824 2704 17888 2706
rect 18112 2704 18176 2706
rect 18400 2704 18464 2706
rect 18688 2704 18752 2706
rect 18976 2704 19040 2706
rect 19264 2704 19328 2706
rect 19552 2704 19616 2706
rect 19840 2704 19904 2706
rect 19978 2698 20054 2706
rect 4282 2622 4358 2630
rect 4714 2622 4790 2630
rect 6154 2622 6230 2630
rect 6586 2622 6662 2630
rect 8746 2622 8822 2630
rect 9754 2622 9830 2630
rect 4282 2620 9830 2622
rect 4282 2564 4292 2620
rect 4348 2564 4724 2620
rect 4780 2564 6164 2620
rect 6220 2564 6596 2620
rect 6652 2564 8756 2620
rect 8812 2564 9764 2620
rect 9820 2564 9830 2620
rect 4282 2562 9830 2564
rect 4282 2554 4358 2562
rect 4714 2554 4790 2562
rect 6154 2554 6230 2562
rect 6586 2554 6662 2562
rect 8746 2554 8822 2562
rect 9754 2554 9830 2562
rect 256 2478 320 2480
rect 826 2478 902 2486
rect 1402 2478 1478 2486
rect 1978 2478 2054 2486
rect 2554 2478 2630 2486
rect 3130 2478 3206 2486
rect 3712 2478 3776 2480
rect 4282 2478 4358 2486
rect 4858 2478 4934 2486
rect 5440 2478 5504 2480
rect 5872 2478 5936 2480
rect 6160 2478 6224 2480
rect 7168 2478 7232 2480
rect 7738 2478 7814 2486
rect 8320 2478 8384 2480
rect 8752 2478 8816 2480
rect 9040 2478 9104 2480
rect 9322 2478 9398 2486
rect 10330 2478 10406 2486
rect 10906 2478 10982 2486
rect 11488 2478 11552 2480
rect 12064 2478 12128 2480
rect 12640 2478 12704 2480
rect 13792 2478 13856 2480
rect 14368 2478 14432 2480
rect 14938 2478 15014 2486
rect 15520 2478 15584 2480
rect 16096 2478 16160 2480
rect 16666 2478 16742 2486
rect 16960 2478 17024 2480
rect 17248 2478 17312 2480
rect 17536 2478 17600 2480
rect 17824 2478 17888 2480
rect 18112 2478 18176 2480
rect 18400 2478 18464 2480
rect 18688 2478 18752 2480
rect 18976 2478 19040 2480
rect 19264 2478 19328 2480
rect 19552 2478 19616 2480
rect 19840 2478 19904 2480
rect 144 2474 432 2478
rect 144 2422 262 2474
rect 314 2422 432 2474
rect 144 2418 432 2422
rect 684 2476 1044 2478
rect 684 2420 836 2476
rect 892 2420 1044 2476
rect 684 2418 1044 2420
rect 1260 2476 1620 2478
rect 1260 2420 1412 2476
rect 1468 2420 1620 2476
rect 1260 2418 1620 2420
rect 1836 2476 2196 2478
rect 1836 2420 1988 2476
rect 2044 2420 2196 2476
rect 1836 2418 2196 2420
rect 2412 2476 2772 2478
rect 2412 2420 2564 2476
rect 2620 2420 2772 2476
rect 2412 2418 2772 2420
rect 2988 2476 3348 2478
rect 2988 2420 3140 2476
rect 3196 2420 3348 2476
rect 2988 2418 3348 2420
rect 3600 2474 3888 2478
rect 3600 2422 3718 2474
rect 3770 2422 3888 2474
rect 3600 2418 3888 2422
rect 4140 2476 4500 2478
rect 4140 2420 4292 2476
rect 4348 2420 4500 2476
rect 4140 2418 4500 2420
rect 4716 2476 5076 2478
rect 4716 2420 4868 2476
rect 4924 2420 5076 2476
rect 4716 2418 5076 2420
rect 5292 2474 6268 2478
rect 5292 2422 5446 2474
rect 5498 2422 5878 2474
rect 5930 2422 6166 2474
rect 6218 2422 6268 2474
rect 5292 2418 6268 2422
rect 7056 2474 7344 2478
rect 7056 2422 7174 2474
rect 7226 2422 7344 2474
rect 7056 2418 7344 2422
rect 7596 2476 7956 2478
rect 7596 2420 7748 2476
rect 7804 2420 7956 2476
rect 7596 2418 7956 2420
rect 8172 2474 9148 2478
rect 8172 2422 8326 2474
rect 8378 2422 8758 2474
rect 8810 2422 9046 2474
rect 9098 2422 9148 2474
rect 8172 2418 9148 2422
rect 9322 2476 10548 2478
rect 9322 2420 9332 2476
rect 9388 2420 10340 2476
rect 10396 2420 10548 2476
rect 9322 2418 10548 2420
rect 10764 2476 11124 2478
rect 10764 2420 10916 2476
rect 10972 2420 11124 2476
rect 10764 2418 11124 2420
rect 11376 2474 11664 2478
rect 11376 2422 11494 2474
rect 11546 2422 11664 2474
rect 11376 2418 11664 2422
rect 11916 2474 12852 2478
rect 11916 2422 12070 2474
rect 12122 2422 12646 2474
rect 12698 2422 12852 2474
rect 11916 2418 12852 2422
rect 13644 2474 14580 2478
rect 13644 2422 13798 2474
rect 13850 2422 14374 2474
rect 14426 2422 14580 2474
rect 13644 2418 14580 2422
rect 14796 2476 15156 2478
rect 14796 2420 14948 2476
rect 15004 2420 15156 2476
rect 14796 2418 15156 2420
rect 15408 2474 15696 2478
rect 15408 2422 15526 2474
rect 15578 2422 15696 2474
rect 15408 2418 15696 2422
rect 15984 2474 16272 2478
rect 15984 2422 16102 2474
rect 16154 2422 16272 2474
rect 15984 2418 16272 2422
rect 16628 2476 19948 2478
rect 16628 2420 16676 2476
rect 16732 2474 19948 2476
rect 16732 2422 16966 2474
rect 17018 2422 17254 2474
rect 17306 2422 17542 2474
rect 17594 2422 17830 2474
rect 17882 2422 18118 2474
rect 18170 2422 18406 2474
rect 18458 2422 18694 2474
rect 18746 2422 18982 2474
rect 19034 2422 19270 2474
rect 19322 2422 19558 2474
rect 19610 2422 19846 2474
rect 19898 2422 19948 2474
rect 16732 2420 19948 2422
rect 16628 2418 19948 2420
rect 256 2416 320 2418
rect 826 2410 902 2418
rect 1402 2410 1478 2418
rect 1978 2410 2054 2418
rect 2554 2410 2630 2418
rect 3130 2410 3206 2418
rect 3712 2416 3776 2418
rect 4282 2410 4358 2418
rect 4858 2410 4934 2418
rect 5440 2416 5504 2418
rect 5872 2416 5936 2418
rect 6160 2416 6224 2418
rect 7168 2416 7232 2418
rect 7738 2410 7814 2418
rect 8320 2416 8384 2418
rect 8752 2416 8816 2418
rect 9040 2416 9104 2418
rect 9322 2410 9398 2418
rect 10330 2410 10406 2418
rect 10906 2410 10982 2418
rect 11488 2416 11552 2418
rect 12064 2416 12128 2418
rect 12640 2416 12704 2418
rect 13792 2416 13856 2418
rect 14368 2416 14432 2418
rect 14938 2410 15014 2418
rect 15520 2416 15584 2418
rect 16096 2416 16160 2418
rect 16666 2410 16742 2418
rect 16960 2416 17024 2418
rect 17248 2416 17312 2418
rect 17536 2416 17600 2418
rect 17824 2416 17888 2418
rect 18112 2416 18176 2418
rect 18400 2416 18464 2418
rect 18688 2416 18752 2418
rect 18976 2416 19040 2418
rect 19264 2416 19328 2418
rect 19552 2416 19616 2418
rect 19840 2416 19904 2418
rect 6010 2334 6086 2342
rect 6730 2334 6806 2342
rect 7594 2334 7670 2342
rect 8890 2334 8966 2342
rect 9610 2334 9686 2342
rect 10186 2334 10262 2342
rect 12496 2334 12560 2336
rect 12784 2334 12848 2336
rect 13648 2334 13712 2336
rect 13930 2334 14006 2342
rect 5868 2332 7670 2334
rect 5868 2276 6020 2332
rect 6076 2276 6740 2332
rect 6796 2276 7604 2332
rect 7660 2276 7670 2332
rect 5868 2274 7670 2276
rect 8748 2332 10262 2334
rect 8748 2276 8900 2332
rect 8956 2276 9620 2332
rect 9676 2276 10196 2332
rect 10252 2276 10262 2332
rect 8748 2274 10262 2276
rect 12452 2332 14044 2334
rect 12452 2330 13940 2332
rect 12452 2278 12502 2330
rect 12554 2278 12790 2330
rect 12842 2278 13654 2330
rect 13706 2278 13940 2330
rect 12452 2276 13940 2278
rect 13996 2276 14044 2332
rect 12452 2274 14044 2276
rect 6010 2266 6086 2274
rect 6730 2266 6806 2274
rect 7594 2266 7670 2274
rect 8890 2266 8966 2274
rect 9610 2266 9686 2274
rect 10186 2266 10262 2274
rect 12496 2272 12560 2274
rect 12784 2272 12848 2274
rect 13648 2272 13712 2274
rect 13930 2266 14006 2274
rect 4858 2190 4934 2198
rect 5866 2190 5942 2198
rect 6874 2190 6950 2198
rect 9034 2190 9110 2198
rect 9466 2190 9542 2198
rect 4858 2188 9542 2190
rect 4858 2132 4868 2188
rect 4924 2132 5876 2188
rect 5932 2132 6884 2188
rect 6940 2132 9044 2188
rect 9100 2132 9476 2188
rect 9532 2132 9542 2188
rect 4858 2130 9542 2132
rect 4858 2122 4934 2130
rect 5866 2122 5942 2130
rect 6874 2122 6950 2130
rect 9034 2122 9110 2130
rect 9466 2122 9542 2130
rect -40 2042 21064 2076
rect -40 1990 118 2042
rect 170 1990 406 2042
rect 458 1990 694 2042
rect 746 1990 982 2042
rect 1034 1990 1270 2042
rect 1322 1990 1558 2042
rect 1610 1990 1846 2042
rect 1898 1990 2134 2042
rect 2186 1990 2422 2042
rect 2474 1990 2710 2042
rect 2762 1990 2998 2042
rect 3050 1990 3286 2042
rect 3338 1990 3574 2042
rect 3626 1990 3862 2042
rect 3914 1990 4150 2042
rect 4202 1990 4438 2042
rect 4490 1990 4726 2042
rect 4778 1990 5014 2042
rect 5066 1990 5302 2042
rect 5354 1990 5590 2042
rect 5642 1990 5878 2042
rect 5930 1990 6166 2042
rect 6218 1990 6454 2042
rect 6506 1990 6742 2042
rect 6794 1990 7030 2042
rect 7082 1990 7318 2042
rect 7370 1990 7606 2042
rect 7658 1990 7894 2042
rect 7946 1990 8182 2042
rect 8234 1990 8470 2042
rect 8522 1990 8758 2042
rect 8810 1990 9046 2042
rect 9098 1990 9334 2042
rect 9386 1990 9622 2042
rect 9674 1990 9910 2042
rect 9962 1990 10198 2042
rect 10250 1990 10486 2042
rect 10538 1990 10774 2042
rect 10826 1990 11062 2042
rect 11114 1990 11350 2042
rect 11402 1990 11638 2042
rect 11690 1990 11926 2042
rect 11978 1990 12214 2042
rect 12266 1990 12502 2042
rect 12554 1990 12790 2042
rect 12842 1990 13078 2042
rect 13130 1990 13366 2042
rect 13418 1990 13654 2042
rect 13706 1990 13942 2042
rect 13994 1990 14230 2042
rect 14282 1990 14518 2042
rect 14570 1990 14806 2042
rect 14858 1990 15094 2042
rect 15146 1990 15382 2042
rect 15434 1990 15670 2042
rect 15722 1990 15958 2042
rect 16010 1990 16246 2042
rect 16298 1990 16534 2042
rect 16586 1990 16822 2042
rect 16874 1990 17110 2042
rect 17162 1990 17398 2042
rect 17450 1990 17686 2042
rect 17738 1990 17974 2042
rect 18026 1990 18262 2042
rect 18314 1990 18550 2042
rect 18602 1990 18838 2042
rect 18890 1990 19126 2042
rect 19178 1990 19414 2042
rect 19466 1990 19702 2042
rect 19754 1990 19990 2042
rect 20042 1990 20278 2042
rect 20330 1990 20566 2042
rect 20618 1990 20854 2042
rect 20906 1990 21064 2042
rect -40 1956 21064 1990
rect 6586 1902 6662 1910
rect 7594 1902 7670 1910
rect 8602 1902 8678 1910
rect 10762 1902 10838 1910
rect 11194 1902 11270 1910
rect 6586 1900 11270 1902
rect 6586 1844 6596 1900
rect 6652 1844 7604 1900
rect 7660 1844 8612 1900
rect 8668 1844 10772 1900
rect 10828 1844 11204 1900
rect 11260 1844 11270 1900
rect 6586 1842 11270 1844
rect 6586 1834 6662 1842
rect 7594 1834 7670 1842
rect 8602 1834 8678 1842
rect 10762 1834 10838 1842
rect 11194 1834 11270 1842
rect 1840 1758 1904 1760
rect 2128 1758 2192 1760
rect 2992 1758 3056 1760
rect 3274 1758 3350 1766
rect 7738 1758 7814 1766
rect 8458 1758 8534 1766
rect 9322 1758 9398 1766
rect 10618 1758 10694 1766
rect 11338 1758 11414 1766
rect 11914 1758 11990 1766
rect 1796 1756 3388 1758
rect 1796 1754 3284 1756
rect 1796 1702 1846 1754
rect 1898 1702 2134 1754
rect 2186 1702 2998 1754
rect 3050 1702 3284 1754
rect 1796 1700 3284 1702
rect 3340 1700 3388 1756
rect 1796 1698 3388 1700
rect 7596 1756 9398 1758
rect 7596 1700 7748 1756
rect 7804 1700 8468 1756
rect 8524 1700 9332 1756
rect 9388 1700 9398 1756
rect 7596 1698 9398 1700
rect 10476 1756 11990 1758
rect 10476 1700 10628 1756
rect 10684 1700 11348 1756
rect 11404 1700 11924 1756
rect 11980 1700 11990 1756
rect 10476 1698 11990 1700
rect 1840 1696 1904 1698
rect 2128 1696 2192 1698
rect 2992 1696 3056 1698
rect 3274 1690 3350 1698
rect 7738 1690 7814 1698
rect 8458 1690 8534 1698
rect 9322 1690 9398 1698
rect 10618 1690 10694 1698
rect 11338 1690 11414 1698
rect 11914 1690 11990 1698
rect 256 1614 320 1616
rect 826 1614 902 1622
rect 1408 1614 1472 1616
rect 1984 1614 2048 1616
rect 3136 1614 3200 1616
rect 3712 1614 3776 1616
rect 4282 1614 4358 1622
rect 4864 1614 4928 1616
rect 5440 1614 5504 1616
rect 6010 1614 6086 1622
rect 6586 1614 6662 1622
rect 7168 1614 7232 1616
rect 7600 1614 7664 1616
rect 7888 1614 7952 1616
rect 8896 1614 8960 1616
rect 9466 1614 9542 1622
rect 10048 1614 10112 1616
rect 10480 1614 10544 1616
rect 10768 1614 10832 1616
rect 11050 1614 11126 1622
rect 12058 1614 12134 1622
rect 12634 1614 12710 1622
rect 13210 1614 13286 1622
rect 13786 1614 13862 1622
rect 14368 1614 14432 1616
rect 14938 1614 15014 1622
rect 15514 1614 15590 1622
rect 16096 1614 16160 1616
rect 16378 1614 16454 1622
rect 16960 1614 17024 1616
rect 17536 1614 17600 1616
rect 17824 1614 17888 1616
rect 18112 1614 18176 1616
rect 18400 1614 18464 1616
rect 18688 1614 18752 1616
rect 18976 1614 19040 1616
rect 19264 1614 19328 1616
rect 19552 1614 19616 1616
rect 19840 1614 19904 1616
rect 20128 1614 20192 1616
rect 20416 1614 20480 1616
rect 20698 1614 20774 1622
rect 144 1610 432 1614
rect 144 1558 262 1610
rect 314 1558 432 1610
rect 144 1554 432 1558
rect 684 1612 1044 1614
rect 684 1556 836 1612
rect 892 1556 1044 1612
rect 684 1554 1044 1556
rect 1260 1610 2196 1614
rect 1260 1558 1414 1610
rect 1466 1558 1990 1610
rect 2042 1558 2196 1610
rect 1260 1554 2196 1558
rect 2988 1610 3924 1614
rect 2988 1558 3142 1610
rect 3194 1558 3718 1610
rect 3770 1558 3924 1610
rect 2988 1554 3924 1558
rect 4140 1612 4500 1614
rect 4140 1556 4292 1612
rect 4348 1556 4500 1612
rect 4140 1554 4500 1556
rect 4752 1610 5040 1614
rect 4752 1558 4870 1610
rect 4922 1558 5040 1610
rect 4752 1554 5040 1558
rect 5328 1610 5616 1614
rect 5328 1558 5446 1610
rect 5498 1558 5616 1610
rect 5328 1554 5616 1558
rect 5868 1612 6228 1614
rect 5868 1556 6020 1612
rect 6076 1556 6228 1612
rect 5868 1554 6228 1556
rect 6444 1612 6804 1614
rect 6444 1556 6596 1612
rect 6652 1556 6804 1612
rect 6444 1554 6804 1556
rect 7020 1610 7996 1614
rect 7020 1558 7174 1610
rect 7226 1558 7606 1610
rect 7658 1558 7894 1610
rect 7946 1558 7996 1610
rect 7020 1554 7996 1558
rect 8784 1610 9072 1614
rect 8784 1558 8902 1610
rect 8954 1558 9072 1610
rect 8784 1554 9072 1558
rect 9324 1612 9684 1614
rect 9324 1556 9476 1612
rect 9532 1556 9684 1612
rect 9324 1554 9684 1556
rect 9900 1610 10876 1614
rect 9900 1558 10054 1610
rect 10106 1558 10486 1610
rect 10538 1558 10774 1610
rect 10826 1558 10876 1610
rect 9900 1554 10876 1558
rect 11050 1612 12276 1614
rect 11050 1556 11060 1612
rect 11116 1556 12068 1612
rect 12124 1556 12276 1612
rect 11050 1554 12276 1556
rect 12492 1612 12852 1614
rect 12492 1556 12644 1612
rect 12700 1556 12852 1612
rect 12492 1554 12852 1556
rect 13068 1612 13428 1614
rect 13068 1556 13220 1612
rect 13276 1556 13428 1612
rect 13068 1554 13428 1556
rect 13644 1612 14004 1614
rect 13644 1556 13796 1612
rect 13852 1556 14004 1612
rect 13644 1554 14004 1556
rect 14256 1610 14544 1614
rect 14256 1558 14374 1610
rect 14426 1558 14544 1610
rect 14256 1554 14544 1558
rect 14796 1612 15156 1614
rect 14796 1556 14948 1612
rect 15004 1556 15156 1612
rect 14796 1554 15156 1556
rect 15372 1612 15732 1614
rect 15372 1556 15524 1612
rect 15580 1556 15732 1612
rect 15372 1554 15732 1556
rect 16052 1612 16492 1614
rect 16052 1610 16388 1612
rect 16052 1558 16102 1610
rect 16154 1558 16388 1610
rect 16052 1556 16388 1558
rect 16444 1556 16492 1612
rect 16052 1554 16492 1556
rect 16848 1610 17136 1614
rect 16848 1558 16966 1610
rect 17018 1558 17136 1610
rect 16848 1554 17136 1558
rect 17492 1612 20812 1614
rect 17492 1610 20708 1612
rect 17492 1558 17542 1610
rect 17594 1558 17830 1610
rect 17882 1558 18118 1610
rect 18170 1558 18406 1610
rect 18458 1558 18694 1610
rect 18746 1558 18982 1610
rect 19034 1558 19270 1610
rect 19322 1558 19558 1610
rect 19610 1558 19846 1610
rect 19898 1558 20134 1610
rect 20186 1558 20422 1610
rect 20474 1558 20708 1610
rect 17492 1556 20708 1558
rect 20764 1556 20812 1612
rect 17492 1554 20812 1556
rect 256 1552 320 1554
rect 826 1546 902 1554
rect 1408 1552 1472 1554
rect 1984 1552 2048 1554
rect 3136 1552 3200 1554
rect 3712 1552 3776 1554
rect 4282 1546 4358 1554
rect 4864 1552 4928 1554
rect 5440 1552 5504 1554
rect 6010 1546 6086 1554
rect 6586 1546 6662 1554
rect 7168 1552 7232 1554
rect 7600 1552 7664 1554
rect 7888 1552 7952 1554
rect 8896 1552 8960 1554
rect 9466 1546 9542 1554
rect 10048 1552 10112 1554
rect 10480 1552 10544 1554
rect 10768 1552 10832 1554
rect 11050 1546 11126 1554
rect 12058 1546 12134 1554
rect 12634 1546 12710 1554
rect 13210 1546 13286 1554
rect 13786 1546 13862 1554
rect 14368 1552 14432 1554
rect 14938 1546 15014 1554
rect 15514 1546 15590 1554
rect 16096 1552 16160 1554
rect 16378 1546 16454 1554
rect 16960 1552 17024 1554
rect 17536 1552 17600 1554
rect 17824 1552 17888 1554
rect 18112 1552 18176 1554
rect 18400 1552 18464 1554
rect 18688 1552 18752 1554
rect 18976 1552 19040 1554
rect 19264 1552 19328 1554
rect 19552 1552 19616 1554
rect 19840 1552 19904 1554
rect 20128 1552 20192 1554
rect 20416 1552 20480 1554
rect 20698 1546 20774 1554
rect 6010 1470 6086 1478
rect 6442 1470 6518 1478
rect 7882 1470 7958 1478
rect 8314 1470 8390 1478
rect 10474 1470 10550 1478
rect 11482 1470 11558 1478
rect 6010 1468 11558 1470
rect 6010 1412 6020 1468
rect 6076 1412 6452 1468
rect 6508 1412 7892 1468
rect 7948 1412 8324 1468
rect 8380 1412 10484 1468
rect 10540 1412 11492 1468
rect 11548 1412 11558 1468
rect 6010 1410 11558 1412
rect 6010 1402 6086 1410
rect 6442 1402 6518 1410
rect 7882 1402 7958 1410
rect 8314 1402 8390 1410
rect 10474 1402 10550 1410
rect 11482 1402 11558 1410
rect 682 1326 758 1334
rect 832 1326 896 1328
rect 1402 1326 1478 1334
rect 1984 1326 2048 1328
rect 2554 1326 2630 1334
rect 682 1324 1044 1326
rect 682 1268 692 1324
rect 748 1322 1044 1324
rect 748 1270 838 1322
rect 890 1270 1044 1322
rect 748 1268 1044 1270
rect 682 1266 1044 1268
rect 1260 1324 1620 1326
rect 1260 1268 1412 1324
rect 1468 1268 1620 1324
rect 1260 1266 1620 1268
rect 1836 1324 2630 1326
rect 1836 1322 2564 1324
rect 1836 1270 1990 1322
rect 2042 1270 2564 1322
rect 1836 1268 2564 1270
rect 2620 1268 2630 1324
rect 1836 1266 2630 1268
rect 682 1258 758 1266
rect 832 1264 896 1266
rect 1402 1258 1478 1266
rect 1984 1264 2048 1266
rect 2554 1258 2630 1266
rect 2842 1326 2918 1334
rect 3136 1326 3200 1328
rect 3706 1326 3782 1334
rect 3994 1326 4070 1334
rect 4288 1326 4352 1328
rect 5866 1326 5942 1334
rect 6016 1326 6080 1328
rect 6442 1326 6518 1334
rect 6592 1326 6656 1328
rect 7162 1326 7238 1334
rect 7744 1326 7808 1328
rect 7882 1326 7958 1334
rect 2842 1324 3348 1326
rect 2842 1268 2852 1324
rect 2908 1322 3348 1324
rect 2908 1270 3142 1322
rect 3194 1270 3348 1322
rect 2908 1268 3348 1270
rect 2842 1266 3348 1268
rect 3564 1324 3924 1326
rect 3564 1268 3716 1324
rect 3772 1268 3924 1324
rect 3564 1266 3924 1268
rect 3994 1324 4500 1326
rect 3994 1268 4004 1324
rect 4060 1322 4500 1324
rect 4060 1270 4294 1322
rect 4346 1270 4500 1322
rect 4060 1268 4500 1270
rect 3994 1266 4500 1268
rect 5866 1324 6228 1326
rect 5866 1268 5876 1324
rect 5932 1322 6228 1324
rect 5932 1270 6022 1322
rect 6074 1270 6228 1322
rect 5932 1268 6228 1270
rect 5866 1266 6228 1268
rect 6442 1324 6804 1326
rect 6442 1268 6452 1324
rect 6508 1322 6804 1324
rect 6508 1270 6598 1322
rect 6650 1270 6804 1322
rect 6508 1268 6804 1270
rect 6442 1266 6804 1268
rect 7020 1324 7380 1326
rect 7020 1268 7172 1324
rect 7228 1268 7380 1324
rect 7020 1266 7380 1268
rect 7596 1324 7958 1326
rect 7596 1322 7892 1324
rect 7596 1270 7750 1322
rect 7802 1270 7892 1322
rect 7596 1268 7892 1270
rect 7948 1268 7958 1324
rect 7596 1266 7958 1268
rect 2842 1258 2918 1266
rect 3136 1264 3200 1266
rect 3706 1258 3782 1266
rect 3994 1258 4070 1266
rect 4288 1264 4352 1266
rect 5866 1258 5942 1266
rect 6016 1264 6080 1266
rect 6442 1258 6518 1266
rect 6592 1264 6656 1266
rect 7162 1258 7238 1266
rect 7744 1264 7808 1266
rect 7882 1258 7958 1266
rect 8464 1326 8528 1328
rect 8602 1326 8678 1334
rect 8464 1324 8678 1326
rect 8464 1322 8612 1324
rect 8464 1270 8470 1322
rect 8522 1270 8612 1322
rect 8464 1268 8612 1270
rect 8668 1268 8678 1324
rect 8464 1266 8678 1268
rect 8464 1264 8528 1266
rect 8602 1258 8678 1266
rect 9322 1326 9398 1334
rect 9472 1326 9536 1328
rect 10042 1326 10118 1334
rect 10624 1326 10688 1328
rect 10762 1326 10838 1334
rect 9322 1324 9684 1326
rect 9322 1268 9332 1324
rect 9388 1322 9684 1324
rect 9388 1270 9478 1322
rect 9530 1270 9684 1322
rect 9388 1268 9684 1270
rect 9322 1266 9684 1268
rect 9900 1324 10260 1326
rect 9900 1268 10052 1324
rect 10108 1268 10260 1324
rect 9900 1266 10260 1268
rect 10476 1324 10838 1326
rect 10476 1322 10772 1324
rect 10476 1270 10630 1322
rect 10682 1270 10772 1322
rect 10476 1268 10772 1270
rect 10828 1268 10838 1324
rect 10476 1266 10838 1268
rect 9322 1258 9398 1266
rect 9472 1264 9536 1266
rect 10042 1258 10118 1266
rect 10624 1264 10688 1266
rect 10762 1258 10838 1266
rect 11344 1326 11408 1328
rect 11482 1326 11558 1334
rect 11344 1324 11558 1326
rect 11344 1322 11492 1324
rect 11344 1270 11350 1322
rect 11402 1270 11492 1322
rect 11344 1268 11492 1270
rect 11548 1268 11558 1324
rect 11344 1266 11558 1268
rect 11344 1264 11408 1266
rect 11482 1258 11558 1266
rect 11914 1326 11990 1334
rect 12064 1326 12128 1328
rect 12490 1326 12566 1334
rect 12640 1326 12704 1328
rect 13066 1326 13142 1334
rect 13216 1326 13280 1328
rect 13642 1326 13718 1334
rect 13792 1326 13856 1328
rect 14794 1326 14870 1334
rect 14944 1326 15008 1328
rect 15520 1326 15584 1328
rect 15658 1326 15734 1334
rect 11914 1324 12276 1326
rect 11914 1268 11924 1324
rect 11980 1322 12276 1324
rect 11980 1270 12070 1322
rect 12122 1270 12276 1322
rect 11980 1268 12276 1270
rect 11914 1266 12276 1268
rect 12490 1324 12852 1326
rect 12490 1268 12500 1324
rect 12556 1322 12852 1324
rect 12556 1270 12646 1322
rect 12698 1270 12852 1322
rect 12556 1268 12852 1270
rect 12490 1266 12852 1268
rect 13066 1324 13428 1326
rect 13066 1268 13076 1324
rect 13132 1322 13428 1324
rect 13132 1270 13222 1322
rect 13274 1270 13428 1322
rect 13132 1268 13428 1270
rect 13066 1266 13428 1268
rect 13642 1324 14004 1326
rect 13642 1268 13652 1324
rect 13708 1322 14004 1324
rect 13708 1270 13798 1322
rect 13850 1270 14004 1322
rect 13708 1268 14004 1270
rect 13642 1266 14004 1268
rect 14794 1324 15156 1326
rect 14794 1268 14804 1324
rect 14860 1322 15156 1324
rect 14860 1270 14950 1322
rect 15002 1270 15156 1322
rect 14860 1268 15156 1270
rect 14794 1266 15156 1268
rect 15372 1324 15734 1326
rect 15372 1322 15668 1324
rect 15372 1270 15526 1322
rect 15578 1270 15668 1322
rect 15372 1268 15668 1270
rect 15724 1268 15734 1324
rect 15372 1266 15734 1268
rect 11914 1258 11990 1266
rect 12064 1264 12128 1266
rect 12490 1258 12566 1266
rect 12640 1264 12704 1266
rect 13066 1258 13142 1266
rect 13216 1264 13280 1266
rect 13642 1258 13718 1266
rect 13792 1264 13856 1266
rect 14794 1258 14870 1266
rect 14944 1264 15008 1266
rect 15520 1264 15584 1266
rect 15658 1258 15734 1266
rect 15946 1326 16022 1334
rect 16096 1326 16160 1328
rect 16384 1326 16448 1328
rect 17386 1326 17462 1334
rect 17536 1326 17600 1328
rect 17824 1326 17888 1328
rect 18112 1326 18176 1328
rect 18400 1326 18464 1328
rect 18688 1326 18752 1328
rect 18976 1326 19040 1328
rect 19264 1326 19328 1328
rect 19552 1326 19616 1328
rect 19840 1326 19904 1328
rect 20128 1326 20192 1328
rect 20416 1326 20480 1328
rect 20704 1326 20768 1328
rect 15946 1324 16492 1326
rect 15946 1268 15956 1324
rect 16012 1322 16492 1324
rect 16012 1270 16102 1322
rect 16154 1270 16390 1322
rect 16442 1270 16492 1322
rect 16012 1268 16492 1270
rect 15946 1266 16492 1268
rect 17386 1324 20812 1326
rect 17386 1268 17396 1324
rect 17452 1322 20812 1324
rect 17452 1270 17542 1322
rect 17594 1270 17830 1322
rect 17882 1270 18118 1322
rect 18170 1270 18406 1322
rect 18458 1270 18694 1322
rect 18746 1270 18982 1322
rect 19034 1270 19270 1322
rect 19322 1270 19558 1322
rect 19610 1270 19846 1322
rect 19898 1270 20134 1322
rect 20186 1270 20422 1322
rect 20474 1270 20710 1322
rect 20762 1270 20812 1322
rect 17452 1268 20812 1270
rect 17386 1266 20812 1268
rect 15946 1258 16022 1266
rect 16096 1264 16160 1266
rect 16384 1264 16448 1266
rect 17386 1258 17462 1266
rect 17536 1264 17600 1266
rect 17824 1264 17888 1266
rect 18112 1264 18176 1266
rect 18400 1264 18464 1266
rect 18688 1264 18752 1266
rect 18976 1264 19040 1266
rect 19264 1264 19328 1266
rect 19552 1264 19616 1266
rect 19840 1264 19904 1266
rect 20128 1264 20192 1266
rect 20416 1264 20480 1266
rect 20704 1264 20768 1266
rect 826 1038 902 1046
rect 2554 1038 2630 1046
rect 826 1036 2630 1038
rect 826 980 836 1036
rect 892 980 2564 1036
rect 2620 980 2630 1036
rect 826 978 2630 980
rect 826 970 902 978
rect 2554 970 2630 978
rect 8170 1038 8246 1046
rect 9466 1038 9542 1046
rect 10042 1038 10118 1046
rect 8170 1036 10118 1038
rect 8170 980 8180 1036
rect 8236 980 9476 1036
rect 9532 980 10052 1036
rect 10108 980 10118 1036
rect 8170 978 10118 980
rect 8170 970 8246 978
rect 9466 970 9542 978
rect 10042 970 10118 978
rect 11050 1038 11126 1046
rect 12634 1038 12710 1046
rect 13066 1038 13142 1046
rect 11050 1036 11396 1038
rect 11050 980 11060 1036
rect 11116 980 11396 1036
rect 11050 978 11396 980
rect 12634 1036 13142 1038
rect 12634 980 12644 1036
rect 12700 980 13076 1036
rect 13132 980 13142 1036
rect 12634 978 13142 980
rect 11050 970 11126 978
rect 12634 970 12710 978
rect 13066 970 13142 978
rect 13786 1038 13862 1046
rect 14794 1038 14870 1046
rect 13786 1036 14870 1038
rect 13786 980 13796 1036
rect 13852 980 14804 1036
rect 14860 980 14870 1036
rect 13786 978 14870 980
rect 13786 970 13862 978
rect 14794 970 14870 978
rect 682 750 758 758
rect 832 750 896 752
rect 1402 750 1478 758
rect 1984 750 2048 752
rect 2266 750 2342 758
rect 682 748 1044 750
rect 682 692 692 748
rect 748 746 1044 748
rect 748 694 838 746
rect 890 694 1044 746
rect 748 692 1044 694
rect 682 690 1044 692
rect 1260 748 1620 750
rect 1260 692 1412 748
rect 1468 692 1620 748
rect 1260 690 1620 692
rect 1836 748 2342 750
rect 1836 746 2276 748
rect 1836 694 1990 746
rect 2042 694 2276 746
rect 1836 692 2276 694
rect 2332 692 2342 748
rect 1836 690 2342 692
rect 682 682 758 690
rect 832 688 896 690
rect 1402 682 1478 690
rect 1984 688 2048 690
rect 2266 682 2342 690
rect 2554 750 2630 758
rect 3136 750 3200 752
rect 3706 750 3782 758
rect 3994 750 4070 758
rect 4288 750 4352 752
rect 5866 750 5942 758
rect 6016 750 6080 752
rect 6442 750 6518 758
rect 6592 750 6656 752
rect 7162 750 7238 758
rect 7594 750 7670 758
rect 7744 750 7808 752
rect 8314 750 8390 758
rect 8464 750 8528 752
rect 2554 748 3348 750
rect 2554 692 2564 748
rect 2620 746 3348 748
rect 2620 694 3142 746
rect 3194 694 3348 746
rect 2620 692 3348 694
rect 2554 690 3348 692
rect 3564 748 3924 750
rect 3564 692 3716 748
rect 3772 692 3924 748
rect 3564 690 3924 692
rect 3994 748 4500 750
rect 3994 692 4004 748
rect 4060 746 4500 748
rect 4060 694 4294 746
rect 4346 694 4500 746
rect 4060 692 4500 694
rect 3994 690 4500 692
rect 5866 748 6228 750
rect 5866 692 5876 748
rect 5932 746 6228 748
rect 5932 694 6022 746
rect 6074 694 6228 746
rect 5932 692 6228 694
rect 5866 690 6228 692
rect 6442 748 6804 750
rect 6442 692 6452 748
rect 6508 746 6804 748
rect 6508 694 6598 746
rect 6650 694 6804 746
rect 6508 692 6804 694
rect 6442 690 6804 692
rect 7020 748 7380 750
rect 7020 692 7172 748
rect 7228 692 7380 748
rect 7020 690 7380 692
rect 7594 748 7956 750
rect 7594 692 7604 748
rect 7660 746 7956 748
rect 7660 694 7750 746
rect 7802 694 7956 746
rect 7660 692 7956 694
rect 7594 690 7956 692
rect 8314 748 8528 750
rect 8314 692 8324 748
rect 8380 746 8528 748
rect 8380 694 8470 746
rect 8522 694 8528 746
rect 8380 692 8528 694
rect 8314 690 8528 692
rect 2554 682 2630 690
rect 3136 688 3200 690
rect 3706 682 3782 690
rect 3994 682 4070 690
rect 4288 688 4352 690
rect 5866 682 5942 690
rect 6016 688 6080 690
rect 6442 682 6518 690
rect 6592 688 6656 690
rect 7162 682 7238 690
rect 7594 682 7670 690
rect 7744 688 7808 690
rect 8314 682 8390 690
rect 8464 688 8528 690
rect 9322 750 9398 758
rect 9472 750 9536 752
rect 10042 750 10118 758
rect 10474 750 10550 758
rect 10624 750 10688 752
rect 11194 750 11270 758
rect 11344 750 11408 752
rect 9322 748 9684 750
rect 9322 692 9332 748
rect 9388 746 9684 748
rect 9388 694 9478 746
rect 9530 694 9684 746
rect 9388 692 9684 694
rect 9322 690 9684 692
rect 9900 748 10260 750
rect 9900 692 10052 748
rect 10108 692 10260 748
rect 9900 690 10260 692
rect 10474 748 10836 750
rect 10474 692 10484 748
rect 10540 746 10836 748
rect 10540 694 10630 746
rect 10682 694 10836 746
rect 10540 692 10836 694
rect 10474 690 10836 692
rect 11194 748 11408 750
rect 11194 692 11204 748
rect 11260 746 11408 748
rect 11260 694 11350 746
rect 11402 694 11408 746
rect 11260 692 11408 694
rect 11194 690 11408 692
rect 9322 682 9398 690
rect 9472 688 9536 690
rect 10042 682 10118 690
rect 10474 682 10550 690
rect 10624 688 10688 690
rect 11194 682 11270 690
rect 11344 688 11408 690
rect 11914 750 11990 758
rect 12064 750 12128 752
rect 12490 750 12566 758
rect 12640 750 12704 752
rect 13066 750 13142 758
rect 13216 750 13280 752
rect 13642 750 13718 758
rect 13792 750 13856 752
rect 14794 750 14870 758
rect 14944 750 15008 752
rect 15520 750 15584 752
rect 15658 750 15734 758
rect 11914 748 12276 750
rect 11914 692 11924 748
rect 11980 746 12276 748
rect 11980 694 12070 746
rect 12122 694 12276 746
rect 11980 692 12276 694
rect 11914 690 12276 692
rect 12490 748 12852 750
rect 12490 692 12500 748
rect 12556 746 12852 748
rect 12556 694 12646 746
rect 12698 694 12852 746
rect 12556 692 12852 694
rect 12490 690 12852 692
rect 13066 748 13428 750
rect 13066 692 13076 748
rect 13132 746 13428 748
rect 13132 694 13222 746
rect 13274 694 13428 746
rect 13132 692 13428 694
rect 13066 690 13428 692
rect 13642 748 14004 750
rect 13642 692 13652 748
rect 13708 746 14004 748
rect 13708 694 13798 746
rect 13850 694 14004 746
rect 13708 692 14004 694
rect 13642 690 14004 692
rect 14794 748 15156 750
rect 14794 692 14804 748
rect 14860 746 15156 748
rect 14860 694 14950 746
rect 15002 694 15156 746
rect 14860 692 15156 694
rect 14794 690 15156 692
rect 15372 748 15734 750
rect 15372 746 15668 748
rect 15372 694 15526 746
rect 15578 694 15668 746
rect 15372 692 15668 694
rect 15724 692 15734 748
rect 15372 690 15734 692
rect 11914 682 11990 690
rect 12064 688 12128 690
rect 12490 682 12566 690
rect 12640 688 12704 690
rect 13066 682 13142 690
rect 13216 688 13280 690
rect 13642 682 13718 690
rect 13792 688 13856 690
rect 14794 682 14870 690
rect 14944 688 15008 690
rect 15520 688 15584 690
rect 15658 682 15734 690
rect 15946 750 16022 758
rect 16096 750 16160 752
rect 16384 750 16448 752
rect 17386 750 17462 758
rect 17536 750 17600 752
rect 17824 750 17888 752
rect 18112 750 18176 752
rect 18400 750 18464 752
rect 18688 750 18752 752
rect 18976 750 19040 752
rect 19264 750 19328 752
rect 19552 750 19616 752
rect 19840 750 19904 752
rect 20128 750 20192 752
rect 20416 750 20480 752
rect 20704 750 20768 752
rect 15946 748 16492 750
rect 15946 692 15956 748
rect 16012 746 16492 748
rect 16012 694 16102 746
rect 16154 694 16390 746
rect 16442 694 16492 746
rect 16012 692 16492 694
rect 15946 690 16492 692
rect 17386 748 20812 750
rect 17386 692 17396 748
rect 17452 746 20812 748
rect 17452 694 17542 746
rect 17594 694 17830 746
rect 17882 694 18118 746
rect 18170 694 18406 746
rect 18458 694 18694 746
rect 18746 694 18982 746
rect 19034 694 19270 746
rect 19322 694 19558 746
rect 19610 694 19846 746
rect 19898 694 20134 746
rect 20186 694 20422 746
rect 20474 694 20710 746
rect 20762 694 20812 746
rect 17452 692 20812 694
rect 17386 690 20812 692
rect 15946 682 16022 690
rect 16096 688 16160 690
rect 16384 688 16448 690
rect 17386 682 17462 690
rect 17536 688 17600 690
rect 17824 688 17888 690
rect 18112 688 18176 690
rect 18400 688 18464 690
rect 18688 688 18752 690
rect 18976 688 19040 690
rect 19264 688 19328 690
rect 19552 688 19616 690
rect 19840 688 19904 690
rect 20128 688 20192 690
rect 20416 688 20480 690
rect 20704 688 20768 690
rect 256 462 320 464
rect 826 462 902 470
rect 1408 462 1472 464
rect 1984 462 2048 464
rect 2266 462 2342 470
rect 2842 462 2918 470
rect 3136 462 3200 464
rect 3712 462 3776 464
rect 4282 462 4358 470
rect 4864 462 4928 464
rect 5440 462 5504 464
rect 6010 462 6086 470
rect 6586 462 6662 470
rect 7168 462 7232 464
rect 7600 462 7664 464
rect 7888 462 7952 464
rect 8896 462 8960 464
rect 9466 462 9542 470
rect 10048 462 10112 464
rect 10480 462 10544 464
rect 10768 462 10832 464
rect 12058 462 12134 470
rect 12634 462 12710 470
rect 13210 462 13286 470
rect 13786 462 13862 470
rect 14368 462 14432 464
rect 14938 462 15014 470
rect 15514 462 15590 470
rect 16096 462 16160 464
rect 16378 462 16454 470
rect 16960 462 17024 464
rect 17536 462 17600 464
rect 17824 462 17888 464
rect 18112 462 18176 464
rect 18400 462 18464 464
rect 18688 462 18752 464
rect 18976 462 19040 464
rect 19264 462 19328 464
rect 19552 462 19616 464
rect 19840 462 19904 464
rect 20128 462 20192 464
rect 20416 462 20480 464
rect 20698 462 20774 470
rect 144 458 432 462
rect 144 406 262 458
rect 314 406 432 458
rect 144 402 432 406
rect 684 460 1044 462
rect 684 404 836 460
rect 892 404 1044 460
rect 684 402 1044 404
rect 1260 458 2196 462
rect 1260 406 1414 458
rect 1466 406 1990 458
rect 2042 406 2196 458
rect 1260 402 2196 406
rect 2266 460 2918 462
rect 2266 404 2276 460
rect 2332 404 2852 460
rect 2908 404 2918 460
rect 2266 402 2918 404
rect 2988 458 3924 462
rect 2988 406 3142 458
rect 3194 406 3718 458
rect 3770 406 3924 458
rect 2988 402 3924 406
rect 4140 460 4500 462
rect 4140 404 4292 460
rect 4348 404 4500 460
rect 4140 402 4500 404
rect 4752 458 5040 462
rect 4752 406 4870 458
rect 4922 406 5040 458
rect 4752 402 5040 406
rect 5328 458 5616 462
rect 5328 406 5446 458
rect 5498 406 5616 458
rect 5328 402 5616 406
rect 5868 460 6228 462
rect 5868 404 6020 460
rect 6076 404 6228 460
rect 5868 402 6228 404
rect 6444 460 6804 462
rect 6444 404 6596 460
rect 6652 404 6804 460
rect 6444 402 6804 404
rect 7020 458 7996 462
rect 7020 406 7174 458
rect 7226 406 7606 458
rect 7658 406 7894 458
rect 7946 406 7996 458
rect 7020 402 7996 406
rect 8784 458 9072 462
rect 8784 406 8902 458
rect 8954 406 9072 458
rect 8784 402 9072 406
rect 9324 460 9684 462
rect 9324 404 9476 460
rect 9532 404 9684 460
rect 9324 402 9684 404
rect 9900 458 10876 462
rect 9900 406 10054 458
rect 10106 406 10486 458
rect 10538 406 10774 458
rect 10826 406 10876 458
rect 9900 402 10876 406
rect 11916 460 12276 462
rect 11916 404 12068 460
rect 12124 404 12276 460
rect 11916 402 12276 404
rect 12492 460 12852 462
rect 12492 404 12644 460
rect 12700 404 12852 460
rect 12492 402 12852 404
rect 13068 460 13428 462
rect 13068 404 13220 460
rect 13276 404 13428 460
rect 13068 402 13428 404
rect 13644 460 14004 462
rect 13644 404 13796 460
rect 13852 404 14004 460
rect 13644 402 14004 404
rect 14256 458 14544 462
rect 14256 406 14374 458
rect 14426 406 14544 458
rect 14256 402 14544 406
rect 14796 460 15156 462
rect 14796 404 14948 460
rect 15004 404 15156 460
rect 14796 402 15156 404
rect 15372 460 15732 462
rect 15372 404 15524 460
rect 15580 404 15732 460
rect 15372 402 15732 404
rect 16052 460 16492 462
rect 16052 458 16388 460
rect 16052 406 16102 458
rect 16154 406 16388 458
rect 16052 404 16388 406
rect 16444 404 16492 460
rect 16052 402 16492 404
rect 16848 458 17136 462
rect 16848 406 16966 458
rect 17018 406 17136 458
rect 16848 402 17136 406
rect 17492 460 20812 462
rect 17492 458 20708 460
rect 17492 406 17542 458
rect 17594 406 17830 458
rect 17882 406 18118 458
rect 18170 406 18406 458
rect 18458 406 18694 458
rect 18746 406 18982 458
rect 19034 406 19270 458
rect 19322 406 19558 458
rect 19610 406 19846 458
rect 19898 406 20134 458
rect 20186 406 20422 458
rect 20474 406 20708 458
rect 17492 404 20708 406
rect 20764 404 20812 460
rect 17492 402 20812 404
rect 256 400 320 402
rect 826 394 902 402
rect 1408 400 1472 402
rect 1984 400 2048 402
rect 2266 394 2342 402
rect 2842 394 2918 402
rect 3136 400 3200 402
rect 3712 400 3776 402
rect 4282 394 4358 402
rect 4864 400 4928 402
rect 5440 400 5504 402
rect 6010 394 6086 402
rect 6586 394 6662 402
rect 7168 400 7232 402
rect 7600 400 7664 402
rect 7888 400 7952 402
rect 8896 400 8960 402
rect 9466 394 9542 402
rect 10048 400 10112 402
rect 10480 400 10544 402
rect 10768 400 10832 402
rect 12058 394 12134 402
rect 12634 394 12710 402
rect 13210 394 13286 402
rect 13786 394 13862 402
rect 14368 400 14432 402
rect 14938 394 15014 402
rect 15514 394 15590 402
rect 16096 400 16160 402
rect 16378 394 16454 402
rect 16960 400 17024 402
rect 17536 400 17600 402
rect 17824 400 17888 402
rect 18112 400 18176 402
rect 18400 400 18464 402
rect 18688 400 18752 402
rect 18976 400 19040 402
rect 19264 400 19328 402
rect 19552 400 19616 402
rect 19840 400 19904 402
rect 20128 400 20192 402
rect 20416 400 20480 402
rect 20698 394 20774 402
rect 1840 318 1904 320
rect 2128 318 2192 320
rect 2992 318 3056 320
rect 3274 318 3350 326
rect 3994 318 4070 326
rect 7738 318 7814 326
rect 1796 316 4070 318
rect 1796 314 3284 316
rect 1796 262 1846 314
rect 1898 262 2134 314
rect 2186 262 2998 314
rect 3050 262 3284 314
rect 1796 260 3284 262
rect 3340 260 4004 316
rect 4060 260 4070 316
rect 1796 258 4070 260
rect 7596 316 7956 318
rect 7596 260 7748 316
rect 7804 260 7956 316
rect 7596 258 7956 260
rect 8458 316 8534 326
rect 10618 318 10694 326
rect 8458 260 8468 316
rect 8524 260 8534 316
rect 1840 256 1904 258
rect 2128 256 2192 258
rect 2992 256 3056 258
rect 3274 250 3350 258
rect 3994 250 4070 258
rect 7738 250 7814 258
rect 8458 250 8534 260
rect 10476 316 10836 318
rect 10476 260 10628 316
rect 10684 260 10836 316
rect 10476 258 10836 260
rect 11338 316 11414 326
rect 11338 260 11348 316
rect 11404 260 11414 316
rect 10618 250 10694 258
rect 11338 250 11414 260
rect -40 26 21064 60
rect -40 -26 118 26
rect 170 -26 406 26
rect 458 -26 694 26
rect 746 -26 982 26
rect 1034 -26 1270 26
rect 1322 -26 1558 26
rect 1610 -26 3574 26
rect 3626 -26 3862 26
rect 3914 -26 4150 26
rect 4202 -26 4438 26
rect 4490 -26 4726 26
rect 4778 -26 5014 26
rect 5066 -26 5302 26
rect 5354 -26 5590 26
rect 5642 -26 5878 26
rect 5930 -26 6166 26
rect 6218 -26 6454 26
rect 6506 -26 6742 26
rect 6794 -26 7030 26
rect 7082 -26 7318 26
rect 7370 -26 8182 26
rect 8234 -26 8758 26
rect 8810 -26 9046 26
rect 9098 -26 9334 26
rect 9386 -26 9622 26
rect 9674 -26 9910 26
rect 9962 -26 10198 26
rect 10250 -26 11062 26
rect 11114 -26 11926 26
rect 11978 -26 12214 26
rect 12266 -26 12502 26
rect 12554 -26 12790 26
rect 12842 -26 13078 26
rect 13130 -26 13366 26
rect 13418 -26 13654 26
rect 13706 -26 13942 26
rect 13994 -26 14230 26
rect 14282 -26 14518 26
rect 14570 -26 14806 26
rect 14858 -26 15094 26
rect 15146 -26 15382 26
rect 15434 -26 15670 26
rect 15722 -26 15958 26
rect 16010 -26 16246 26
rect 16298 -26 16534 26
rect 16586 -26 16822 26
rect 16874 -26 17110 26
rect 17162 -26 17398 26
rect 17450 -26 17686 26
rect 17738 -26 17974 26
rect 18026 -26 18262 26
rect 18314 -26 18550 26
rect 18602 -26 18838 26
rect 18890 -26 19126 26
rect 19178 -26 19414 26
rect 19466 -26 19702 26
rect 19754 -26 19990 26
rect 20042 -26 20278 26
rect 20330 -26 20566 26
rect 20618 -26 20854 26
rect 20906 -26 21064 26
rect -40 -60 21064 -26
<< via2 >>
rect 6020 3770 6076 3772
rect 6020 3718 6022 3770
rect 6022 3718 6074 3770
rect 6074 3718 6076 3770
rect 6020 3716 6076 3718
rect 6740 3770 6796 3772
rect 6740 3718 6742 3770
rect 6742 3718 6794 3770
rect 6794 3718 6796 3770
rect 6740 3716 6796 3718
rect 8900 3770 8956 3772
rect 8900 3718 8902 3770
rect 8902 3718 8954 3770
rect 8954 3718 8956 3770
rect 8900 3716 8956 3718
rect 9620 3770 9676 3772
rect 9620 3718 9622 3770
rect 9622 3718 9674 3770
rect 9674 3718 9676 3770
rect 9620 3716 9676 3718
rect 13940 3770 13996 3772
rect 13940 3718 13942 3770
rect 13942 3718 13994 3770
rect 13994 3718 13996 3770
rect 13940 3716 13996 3718
rect 14660 3716 14716 3772
rect 836 3626 892 3628
rect 836 3574 838 3626
rect 838 3574 890 3626
rect 890 3574 892 3626
rect 836 3572 892 3574
rect 1412 3626 1468 3628
rect 1412 3574 1414 3626
rect 1414 3574 1466 3626
rect 1466 3574 1468 3626
rect 1412 3572 1468 3574
rect 1988 3626 2044 3628
rect 1988 3574 1990 3626
rect 1990 3574 2042 3626
rect 2042 3574 2044 3626
rect 1988 3572 2044 3574
rect 2564 3626 2620 3628
rect 2564 3574 2566 3626
rect 2566 3574 2618 3626
rect 2618 3574 2620 3626
rect 2564 3572 2620 3574
rect 3140 3626 3196 3628
rect 3140 3574 3142 3626
rect 3142 3574 3194 3626
rect 3194 3574 3196 3626
rect 3140 3572 3196 3574
rect 4292 3626 4348 3628
rect 4292 3574 4294 3626
rect 4294 3574 4346 3626
rect 4346 3574 4348 3626
rect 4292 3572 4348 3574
rect 4868 3626 4924 3628
rect 4868 3574 4870 3626
rect 4870 3574 4922 3626
rect 4922 3574 4924 3626
rect 4868 3572 4924 3574
rect 7748 3626 7804 3628
rect 7748 3574 7750 3626
rect 7750 3574 7802 3626
rect 7802 3574 7804 3626
rect 7748 3572 7804 3574
rect 10340 3626 10396 3628
rect 10340 3574 10342 3626
rect 10342 3574 10394 3626
rect 10394 3574 10396 3626
rect 10340 3572 10396 3574
rect 10916 3626 10972 3628
rect 10916 3574 10918 3626
rect 10918 3574 10970 3626
rect 10970 3574 10972 3626
rect 10916 3572 10972 3574
rect 12932 3572 12988 3628
rect 13508 3572 13564 3628
rect 14948 3626 15004 3628
rect 14948 3574 14950 3626
rect 14950 3574 15002 3626
rect 15002 3574 15004 3626
rect 14948 3572 15004 3574
rect 16676 3626 16732 3628
rect 16676 3574 16678 3626
rect 16678 3574 16730 3626
rect 16730 3574 16732 3626
rect 16676 3572 16732 3574
rect 980 3284 1036 3340
rect 1556 3284 1612 3340
rect 2132 3284 2188 3340
rect 2708 3284 2764 3340
rect 2996 3284 3052 3340
rect 4148 3284 4204 3340
rect 4724 3284 4780 3340
rect 5444 3338 5500 3340
rect 5444 3286 5446 3338
rect 5446 3286 5498 3338
rect 5498 3286 5500 3338
rect 5444 3284 5500 3286
rect 5876 3284 5932 3340
rect 6596 3284 6652 3340
rect 7604 3284 7660 3340
rect 8324 3338 8380 3340
rect 8324 3286 8326 3338
rect 8326 3286 8378 3338
rect 8378 3286 8380 3338
rect 8324 3284 8380 3286
rect 8756 3284 8812 3340
rect 9476 3284 9532 3340
rect 10196 3284 10252 3340
rect 10772 3284 10828 3340
rect 12068 3338 12124 3340
rect 12068 3286 12070 3338
rect 12070 3286 12122 3338
rect 12122 3286 12124 3338
rect 12068 3284 12124 3286
rect 12932 3284 12988 3340
rect 13220 3284 13276 3340
rect 14372 3338 14428 3340
rect 14372 3286 14374 3338
rect 14374 3286 14426 3338
rect 14426 3286 14428 3338
rect 14372 3284 14428 3286
rect 14660 3284 14716 3340
rect 19988 3284 20044 3340
rect 1556 2996 1612 3052
rect 1988 2996 2044 3052
rect 6452 3050 6508 3052
rect 6452 2998 6454 3050
rect 6454 2998 6506 3050
rect 6506 2998 6508 3050
rect 6452 2996 6508 2998
rect 7748 2996 7804 3052
rect 8324 2996 8380 3052
rect 9332 3050 9388 3052
rect 9332 2998 9334 3050
rect 9334 2998 9386 3050
rect 9386 2998 9388 3050
rect 9332 2996 9388 2998
rect 980 2708 1036 2764
rect 1556 2708 1612 2764
rect 2132 2708 2188 2764
rect 2708 2708 2764 2764
rect 2996 2708 3052 2764
rect 4148 2708 4204 2764
rect 4724 2708 4780 2764
rect 5444 2762 5500 2764
rect 5444 2710 5446 2762
rect 5446 2710 5498 2762
rect 5498 2710 5500 2762
rect 5444 2708 5500 2710
rect 6164 2708 6220 2764
rect 6884 2708 6940 2764
rect 7604 2708 7660 2764
rect 8324 2762 8380 2764
rect 8324 2710 8326 2762
rect 8326 2710 8378 2762
rect 8378 2710 8380 2762
rect 8324 2708 8380 2710
rect 9044 2708 9100 2764
rect 9764 2708 9820 2764
rect 10196 2708 10252 2764
rect 10772 2708 10828 2764
rect 12068 2762 12124 2764
rect 12068 2710 12070 2762
rect 12070 2710 12122 2762
rect 12122 2710 12124 2762
rect 12068 2708 12124 2710
rect 13220 2708 13276 2764
rect 13508 2708 13564 2764
rect 14372 2762 14428 2764
rect 14372 2710 14374 2762
rect 14374 2710 14426 2762
rect 14426 2710 14428 2762
rect 14372 2708 14428 2710
rect 14660 2708 14716 2764
rect 19988 2708 20044 2764
rect 4292 2564 4348 2620
rect 4724 2564 4780 2620
rect 6164 2564 6220 2620
rect 6596 2564 6652 2620
rect 8756 2564 8812 2620
rect 9764 2564 9820 2620
rect 836 2474 892 2476
rect 836 2422 838 2474
rect 838 2422 890 2474
rect 890 2422 892 2474
rect 836 2420 892 2422
rect 1412 2474 1468 2476
rect 1412 2422 1414 2474
rect 1414 2422 1466 2474
rect 1466 2422 1468 2474
rect 1412 2420 1468 2422
rect 1988 2474 2044 2476
rect 1988 2422 1990 2474
rect 1990 2422 2042 2474
rect 2042 2422 2044 2474
rect 1988 2420 2044 2422
rect 2564 2474 2620 2476
rect 2564 2422 2566 2474
rect 2566 2422 2618 2474
rect 2618 2422 2620 2474
rect 2564 2420 2620 2422
rect 3140 2474 3196 2476
rect 3140 2422 3142 2474
rect 3142 2422 3194 2474
rect 3194 2422 3196 2474
rect 3140 2420 3196 2422
rect 4292 2474 4348 2476
rect 4292 2422 4294 2474
rect 4294 2422 4346 2474
rect 4346 2422 4348 2474
rect 4292 2420 4348 2422
rect 4868 2474 4924 2476
rect 4868 2422 4870 2474
rect 4870 2422 4922 2474
rect 4922 2422 4924 2474
rect 4868 2420 4924 2422
rect 7748 2474 7804 2476
rect 7748 2422 7750 2474
rect 7750 2422 7802 2474
rect 7802 2422 7804 2474
rect 7748 2420 7804 2422
rect 9332 2420 9388 2476
rect 10340 2474 10396 2476
rect 10340 2422 10342 2474
rect 10342 2422 10394 2474
rect 10394 2422 10396 2474
rect 10340 2420 10396 2422
rect 10916 2474 10972 2476
rect 10916 2422 10918 2474
rect 10918 2422 10970 2474
rect 10970 2422 10972 2474
rect 10916 2420 10972 2422
rect 14948 2474 15004 2476
rect 14948 2422 14950 2474
rect 14950 2422 15002 2474
rect 15002 2422 15004 2474
rect 14948 2420 15004 2422
rect 16676 2474 16732 2476
rect 16676 2422 16678 2474
rect 16678 2422 16730 2474
rect 16730 2422 16732 2474
rect 16676 2420 16732 2422
rect 6020 2330 6076 2332
rect 6020 2278 6022 2330
rect 6022 2278 6074 2330
rect 6074 2278 6076 2330
rect 6020 2276 6076 2278
rect 6740 2330 6796 2332
rect 6740 2278 6742 2330
rect 6742 2278 6794 2330
rect 6794 2278 6796 2330
rect 6740 2276 6796 2278
rect 7604 2276 7660 2332
rect 8900 2330 8956 2332
rect 8900 2278 8902 2330
rect 8902 2278 8954 2330
rect 8954 2278 8956 2330
rect 8900 2276 8956 2278
rect 9620 2330 9676 2332
rect 9620 2278 9622 2330
rect 9622 2278 9674 2330
rect 9674 2278 9676 2330
rect 9620 2276 9676 2278
rect 10196 2276 10252 2332
rect 13940 2330 13996 2332
rect 13940 2278 13942 2330
rect 13942 2278 13994 2330
rect 13994 2278 13996 2330
rect 13940 2276 13996 2278
rect 4868 2132 4924 2188
rect 5876 2132 5932 2188
rect 6884 2132 6940 2188
rect 9044 2132 9100 2188
rect 9476 2132 9532 2188
rect 6596 1844 6652 1900
rect 7604 1844 7660 1900
rect 8612 1844 8668 1900
rect 10772 1844 10828 1900
rect 11204 1844 11260 1900
rect 3284 1754 3340 1756
rect 3284 1702 3286 1754
rect 3286 1702 3338 1754
rect 3338 1702 3340 1754
rect 3284 1700 3340 1702
rect 7748 1754 7804 1756
rect 7748 1702 7750 1754
rect 7750 1702 7802 1754
rect 7802 1702 7804 1754
rect 7748 1700 7804 1702
rect 8468 1754 8524 1756
rect 8468 1702 8470 1754
rect 8470 1702 8522 1754
rect 8522 1702 8524 1754
rect 8468 1700 8524 1702
rect 9332 1700 9388 1756
rect 10628 1754 10684 1756
rect 10628 1702 10630 1754
rect 10630 1702 10682 1754
rect 10682 1702 10684 1754
rect 10628 1700 10684 1702
rect 11348 1754 11404 1756
rect 11348 1702 11350 1754
rect 11350 1702 11402 1754
rect 11402 1702 11404 1754
rect 11348 1700 11404 1702
rect 11924 1700 11980 1756
rect 836 1610 892 1612
rect 836 1558 838 1610
rect 838 1558 890 1610
rect 890 1558 892 1610
rect 836 1556 892 1558
rect 4292 1610 4348 1612
rect 4292 1558 4294 1610
rect 4294 1558 4346 1610
rect 4346 1558 4348 1610
rect 4292 1556 4348 1558
rect 6020 1610 6076 1612
rect 6020 1558 6022 1610
rect 6022 1558 6074 1610
rect 6074 1558 6076 1610
rect 6020 1556 6076 1558
rect 6596 1610 6652 1612
rect 6596 1558 6598 1610
rect 6598 1558 6650 1610
rect 6650 1558 6652 1610
rect 6596 1556 6652 1558
rect 9476 1610 9532 1612
rect 9476 1558 9478 1610
rect 9478 1558 9530 1610
rect 9530 1558 9532 1610
rect 9476 1556 9532 1558
rect 11060 1556 11116 1612
rect 12068 1610 12124 1612
rect 12068 1558 12070 1610
rect 12070 1558 12122 1610
rect 12122 1558 12124 1610
rect 12068 1556 12124 1558
rect 12644 1610 12700 1612
rect 12644 1558 12646 1610
rect 12646 1558 12698 1610
rect 12698 1558 12700 1610
rect 12644 1556 12700 1558
rect 13220 1610 13276 1612
rect 13220 1558 13222 1610
rect 13222 1558 13274 1610
rect 13274 1558 13276 1610
rect 13220 1556 13276 1558
rect 13796 1610 13852 1612
rect 13796 1558 13798 1610
rect 13798 1558 13850 1610
rect 13850 1558 13852 1610
rect 13796 1556 13852 1558
rect 14948 1610 15004 1612
rect 14948 1558 14950 1610
rect 14950 1558 15002 1610
rect 15002 1558 15004 1610
rect 14948 1556 15004 1558
rect 15524 1610 15580 1612
rect 15524 1558 15526 1610
rect 15526 1558 15578 1610
rect 15578 1558 15580 1610
rect 15524 1556 15580 1558
rect 16388 1610 16444 1612
rect 16388 1558 16390 1610
rect 16390 1558 16442 1610
rect 16442 1558 16444 1610
rect 16388 1556 16444 1558
rect 20708 1610 20764 1612
rect 20708 1558 20710 1610
rect 20710 1558 20762 1610
rect 20762 1558 20764 1610
rect 20708 1556 20764 1558
rect 6020 1412 6076 1468
rect 6452 1412 6508 1468
rect 7892 1412 7948 1468
rect 8324 1412 8380 1468
rect 10484 1412 10540 1468
rect 11492 1412 11548 1468
rect 692 1268 748 1324
rect 1412 1322 1468 1324
rect 1412 1270 1414 1322
rect 1414 1270 1466 1322
rect 1466 1270 1468 1322
rect 1412 1268 1468 1270
rect 2564 1268 2620 1324
rect 2852 1268 2908 1324
rect 3716 1322 3772 1324
rect 3716 1270 3718 1322
rect 3718 1270 3770 1322
rect 3770 1270 3772 1322
rect 3716 1268 3772 1270
rect 4004 1268 4060 1324
rect 5876 1268 5932 1324
rect 6452 1268 6508 1324
rect 7172 1322 7228 1324
rect 7172 1270 7174 1322
rect 7174 1270 7226 1322
rect 7226 1270 7228 1322
rect 7172 1268 7228 1270
rect 7892 1268 7948 1324
rect 8612 1268 8668 1324
rect 9332 1268 9388 1324
rect 10052 1322 10108 1324
rect 10052 1270 10054 1322
rect 10054 1270 10106 1322
rect 10106 1270 10108 1322
rect 10052 1268 10108 1270
rect 10772 1268 10828 1324
rect 11492 1268 11548 1324
rect 11924 1268 11980 1324
rect 12500 1268 12556 1324
rect 13076 1268 13132 1324
rect 13652 1268 13708 1324
rect 14804 1268 14860 1324
rect 15668 1268 15724 1324
rect 15956 1268 16012 1324
rect 17396 1268 17452 1324
rect 836 980 892 1036
rect 2564 980 2620 1036
rect 8180 1034 8236 1036
rect 8180 982 8182 1034
rect 8182 982 8234 1034
rect 8234 982 8236 1034
rect 8180 980 8236 982
rect 9476 980 9532 1036
rect 10052 980 10108 1036
rect 11060 1034 11116 1036
rect 11060 982 11062 1034
rect 11062 982 11114 1034
rect 11114 982 11116 1034
rect 11060 980 11116 982
rect 12644 980 12700 1036
rect 13076 980 13132 1036
rect 13796 980 13852 1036
rect 14804 980 14860 1036
rect 692 692 748 748
rect 1412 746 1468 748
rect 1412 694 1414 746
rect 1414 694 1466 746
rect 1466 694 1468 746
rect 1412 692 1468 694
rect 2276 692 2332 748
rect 2564 692 2620 748
rect 3716 746 3772 748
rect 3716 694 3718 746
rect 3718 694 3770 746
rect 3770 694 3772 746
rect 3716 692 3772 694
rect 4004 692 4060 748
rect 5876 692 5932 748
rect 6452 692 6508 748
rect 7172 746 7228 748
rect 7172 694 7174 746
rect 7174 694 7226 746
rect 7226 694 7228 746
rect 7172 692 7228 694
rect 7604 692 7660 748
rect 8324 692 8380 748
rect 9332 692 9388 748
rect 10052 746 10108 748
rect 10052 694 10054 746
rect 10054 694 10106 746
rect 10106 694 10108 746
rect 10052 692 10108 694
rect 10484 692 10540 748
rect 11204 692 11260 748
rect 11924 692 11980 748
rect 12500 692 12556 748
rect 13076 692 13132 748
rect 13652 692 13708 748
rect 14804 692 14860 748
rect 15668 692 15724 748
rect 15956 692 16012 748
rect 17396 692 17452 748
rect 836 458 892 460
rect 836 406 838 458
rect 838 406 890 458
rect 890 406 892 458
rect 836 404 892 406
rect 2276 404 2332 460
rect 2852 404 2908 460
rect 4292 458 4348 460
rect 4292 406 4294 458
rect 4294 406 4346 458
rect 4346 406 4348 458
rect 4292 404 4348 406
rect 6020 458 6076 460
rect 6020 406 6022 458
rect 6022 406 6074 458
rect 6074 406 6076 458
rect 6020 404 6076 406
rect 6596 458 6652 460
rect 6596 406 6598 458
rect 6598 406 6650 458
rect 6650 406 6652 458
rect 6596 404 6652 406
rect 9476 458 9532 460
rect 9476 406 9478 458
rect 9478 406 9530 458
rect 9530 406 9532 458
rect 9476 404 9532 406
rect 12068 458 12124 460
rect 12068 406 12070 458
rect 12070 406 12122 458
rect 12122 406 12124 458
rect 12068 404 12124 406
rect 12644 458 12700 460
rect 12644 406 12646 458
rect 12646 406 12698 458
rect 12698 406 12700 458
rect 12644 404 12700 406
rect 13220 458 13276 460
rect 13220 406 13222 458
rect 13222 406 13274 458
rect 13274 406 13276 458
rect 13220 404 13276 406
rect 13796 458 13852 460
rect 13796 406 13798 458
rect 13798 406 13850 458
rect 13850 406 13852 458
rect 13796 404 13852 406
rect 14948 458 15004 460
rect 14948 406 14950 458
rect 14950 406 15002 458
rect 15002 406 15004 458
rect 14948 404 15004 406
rect 15524 458 15580 460
rect 15524 406 15526 458
rect 15526 406 15578 458
rect 15578 406 15580 458
rect 15524 404 15580 406
rect 16388 458 16444 460
rect 16388 406 16390 458
rect 16390 406 16442 458
rect 16442 406 16444 458
rect 16388 404 16444 406
rect 20708 458 20764 460
rect 20708 406 20710 458
rect 20710 406 20762 458
rect 20762 406 20764 458
rect 20708 404 20764 406
rect 3284 314 3340 316
rect 3284 262 3286 314
rect 3286 262 3338 314
rect 3338 262 3340 314
rect 3284 260 3340 262
rect 4004 260 4060 316
rect 7748 314 7804 316
rect 7748 262 7750 314
rect 7750 262 7802 314
rect 7802 262 7804 314
rect 7748 260 7804 262
rect 8468 314 8524 316
rect 8468 262 8470 314
rect 8470 262 8522 314
rect 8522 262 8524 314
rect 8468 260 8524 262
rect 10628 314 10684 316
rect 10628 262 10630 314
rect 10630 262 10682 314
rect 10682 262 10684 314
rect 10628 260 10684 262
rect 11348 314 11404 316
rect 11348 262 11350 314
rect 11350 262 11402 314
rect 11402 262 11404 314
rect 11348 260 11404 262
<< metal3 >>
rect 6010 3772 6086 3782
rect 6010 3716 6020 3772
rect 6076 3716 6086 3772
rect 6010 3706 6086 3716
rect 6730 3772 6806 3782
rect 6730 3716 6740 3772
rect 6796 3716 6806 3772
rect 6730 3706 6806 3716
rect 8890 3772 8966 3782
rect 8890 3716 8900 3772
rect 8956 3716 8966 3772
rect 8890 3706 8966 3716
rect 9610 3772 9686 3782
rect 9610 3716 9620 3772
rect 9676 3716 9686 3772
rect 9610 3706 9686 3716
rect 826 3628 902 3638
rect 826 3572 836 3628
rect 892 3572 902 3628
rect 826 3562 902 3572
rect 1402 3628 1478 3638
rect 1402 3572 1412 3628
rect 1468 3572 1478 3628
rect 1402 3562 1478 3572
rect 1978 3628 2054 3638
rect 1978 3572 1988 3628
rect 2044 3572 2054 3628
rect 1978 3562 2054 3572
rect 2554 3628 2630 3638
rect 2554 3572 2564 3628
rect 2620 3572 2630 3628
rect 2554 3562 2630 3572
rect 3130 3628 3206 3638
rect 3130 3572 3140 3628
rect 3196 3572 3206 3628
rect 3130 3562 3206 3572
rect 4282 3628 4358 3638
rect 4282 3572 4292 3628
rect 4348 3572 4358 3628
rect 4282 3562 4358 3572
rect 4858 3628 4934 3638
rect 4858 3572 4868 3628
rect 4924 3572 4934 3628
rect 4858 3562 4934 3572
rect 834 2486 894 3562
rect 970 3340 1046 3350
rect 970 3284 980 3340
rect 1036 3284 1046 3340
rect 970 3274 1046 3284
rect 978 2774 1038 3274
rect 1410 2774 1470 3562
rect 1546 3340 1622 3350
rect 1546 3284 1556 3340
rect 1612 3284 1622 3340
rect 1546 3274 1622 3284
rect 1554 3062 1614 3274
rect 1986 3062 2046 3562
rect 2122 3340 2198 3350
rect 2122 3284 2132 3340
rect 2188 3284 2198 3340
rect 2122 3274 2198 3284
rect 1546 3052 1622 3062
rect 1546 2996 1556 3052
rect 1612 2996 1622 3052
rect 1546 2986 1622 2996
rect 1978 3052 2054 3062
rect 1978 2996 1988 3052
rect 2044 2996 2054 3052
rect 1978 2986 2054 2996
rect 1554 2774 1614 2986
rect 970 2768 1046 2774
rect 970 2704 976 2768
rect 1040 2704 1046 2768
rect 970 2698 1046 2704
rect 1402 2768 1478 2774
rect 1402 2704 1408 2768
rect 1472 2704 1478 2768
rect 1402 2698 1478 2704
rect 1546 2764 1622 2774
rect 1546 2708 1556 2764
rect 1612 2708 1622 2764
rect 1546 2698 1622 2708
rect 1410 2486 1470 2698
rect 1986 2486 2046 2986
rect 2130 2774 2190 3274
rect 2562 2774 2622 3562
rect 2698 3340 2774 3350
rect 2698 3284 2708 3340
rect 2764 3284 2774 3340
rect 2698 3274 2774 3284
rect 2986 3340 3062 3350
rect 2986 3284 2996 3340
rect 3052 3284 3062 3340
rect 2986 3274 3062 3284
rect 2706 2774 2766 3274
rect 2994 2774 3054 3274
rect 3138 2774 3198 3562
rect 4138 3340 4214 3350
rect 4138 3284 4148 3340
rect 4204 3284 4214 3340
rect 4138 3274 4214 3284
rect 4146 2774 4206 3274
rect 2122 2768 2198 2774
rect 2122 2704 2128 2768
rect 2192 2704 2198 2768
rect 2122 2698 2198 2704
rect 2554 2768 2630 2774
rect 2554 2704 2560 2768
rect 2624 2704 2630 2768
rect 2554 2698 2630 2704
rect 2698 2764 2774 2774
rect 2698 2708 2708 2764
rect 2764 2708 2774 2764
rect 2698 2698 2774 2708
rect 2986 2764 3062 2774
rect 2986 2708 2996 2764
rect 3052 2708 3062 2764
rect 2986 2698 3062 2708
rect 3130 2768 3206 2774
rect 3130 2704 3136 2768
rect 3200 2704 3206 2768
rect 3130 2698 3206 2704
rect 4138 2768 4214 2774
rect 4138 2704 4144 2768
rect 4208 2704 4214 2768
rect 4138 2698 4214 2704
rect 2562 2486 2622 2698
rect 826 2476 902 2486
rect 826 2420 836 2476
rect 892 2420 902 2476
rect 826 2410 902 2420
rect 1402 2476 1478 2486
rect 1402 2420 1412 2476
rect 1468 2420 1478 2476
rect 1402 2410 1478 2420
rect 1978 2476 2054 2486
rect 1978 2420 1988 2476
rect 2044 2420 2054 2476
rect 1978 2410 2054 2420
rect 2554 2476 2630 2486
rect 2554 2420 2564 2476
rect 2620 2420 2630 2476
rect 2554 2410 2630 2420
rect 2706 1910 2766 2698
rect 3138 2486 3198 2698
rect 4290 2630 4350 3562
rect 4714 3340 4790 3350
rect 4714 3284 4724 3340
rect 4780 3284 4790 3340
rect 4714 3274 4790 3284
rect 4722 2774 4782 3274
rect 4714 2764 4790 2774
rect 4714 2708 4724 2764
rect 4780 2708 4790 2764
rect 4714 2698 4790 2708
rect 4722 2630 4782 2698
rect 4282 2620 4358 2630
rect 4282 2564 4292 2620
rect 4348 2564 4358 2620
rect 4282 2554 4358 2564
rect 4714 2620 4790 2630
rect 4714 2564 4724 2620
rect 4780 2564 4790 2620
rect 4714 2554 4790 2564
rect 4290 2486 4350 2554
rect 4866 2486 4926 3562
rect 5434 3340 5510 3350
rect 5434 3284 5444 3340
rect 5500 3284 5510 3340
rect 5434 3274 5510 3284
rect 5866 3340 5942 3350
rect 5866 3284 5876 3340
rect 5932 3284 5942 3340
rect 5866 3274 5942 3284
rect 5442 2774 5502 3274
rect 5434 2768 5510 2774
rect 5434 2704 5440 2768
rect 5504 2704 5510 2768
rect 5434 2698 5510 2704
rect 3130 2476 3206 2486
rect 3130 2420 3140 2476
rect 3196 2420 3206 2476
rect 3130 2410 3206 2420
rect 4282 2476 4358 2486
rect 4282 2420 4292 2476
rect 4348 2420 4358 2476
rect 4282 2410 4358 2420
rect 4858 2476 4934 2486
rect 4858 2420 4868 2476
rect 4924 2420 4934 2476
rect 4858 2410 4934 2420
rect 4866 2198 4926 2410
rect 5874 2198 5934 3274
rect 6018 2342 6078 3706
rect 6162 2774 6222 3342
rect 6450 3062 6510 3342
rect 6586 3340 6662 3350
rect 6586 3284 6596 3340
rect 6652 3284 6662 3340
rect 6586 3274 6662 3284
rect 6442 3052 6518 3062
rect 6442 2996 6452 3052
rect 6508 2996 6518 3052
rect 6442 2986 6518 2996
rect 6154 2764 6230 2774
rect 6154 2708 6164 2764
rect 6220 2708 6230 2764
rect 6154 2698 6230 2708
rect 6450 2706 6510 2986
rect 6162 2630 6222 2698
rect 6594 2630 6654 3274
rect 6154 2620 6230 2630
rect 6154 2564 6164 2620
rect 6220 2564 6230 2620
rect 6154 2554 6230 2564
rect 6586 2620 6662 2630
rect 6586 2564 6596 2620
rect 6652 2564 6662 2620
rect 6586 2554 6662 2564
rect 6738 2342 6798 3706
rect 7738 3628 7814 3638
rect 7738 3572 7748 3628
rect 7804 3572 7814 3628
rect 7738 3562 7814 3572
rect 6882 2774 6942 3342
rect 7594 3340 7670 3350
rect 7594 3284 7604 3340
rect 7660 3284 7670 3340
rect 7594 3274 7670 3284
rect 7602 2774 7662 3274
rect 7746 3062 7806 3562
rect 8314 3340 8390 3350
rect 8314 3284 8324 3340
rect 8380 3284 8390 3340
rect 8314 3274 8390 3284
rect 8746 3340 8822 3350
rect 8746 3284 8756 3340
rect 8812 3284 8822 3340
rect 8746 3274 8822 3284
rect 8322 3062 8382 3274
rect 7738 3052 7814 3062
rect 7738 2996 7748 3052
rect 7804 2996 7814 3052
rect 7738 2986 7814 2996
rect 8314 3052 8390 3062
rect 8314 2996 8324 3052
rect 8380 2996 8390 3052
rect 8314 2986 8390 2996
rect 6874 2764 6950 2774
rect 6874 2708 6884 2764
rect 6940 2708 6950 2764
rect 6874 2698 6950 2708
rect 7594 2764 7670 2774
rect 7594 2708 7604 2764
rect 7660 2708 7670 2764
rect 7594 2698 7670 2708
rect 6010 2332 6086 2342
rect 6010 2276 6020 2332
rect 6076 2276 6086 2332
rect 6010 2266 6086 2276
rect 6730 2332 6806 2342
rect 6730 2276 6740 2332
rect 6796 2276 6806 2332
rect 6730 2266 6806 2276
rect 6882 2198 6942 2698
rect 7602 2342 7662 2698
rect 7746 2486 7806 2986
rect 8322 2774 8382 2986
rect 8314 2764 8390 2774
rect 8314 2708 8324 2764
rect 8380 2708 8390 2764
rect 8314 2698 8390 2708
rect 8754 2630 8814 3274
rect 8746 2620 8822 2630
rect 8746 2564 8756 2620
rect 8812 2564 8822 2620
rect 8746 2554 8822 2564
rect 7738 2476 7814 2486
rect 7738 2420 7748 2476
rect 7804 2420 7814 2476
rect 7738 2410 7814 2420
rect 8898 2342 8958 3706
rect 9042 2774 9102 3342
rect 9330 3062 9390 3342
rect 9466 3340 9542 3350
rect 9466 3284 9476 3340
rect 9532 3284 9542 3340
rect 9466 3274 9542 3284
rect 9322 3052 9398 3062
rect 9322 2996 9332 3052
rect 9388 2996 9398 3052
rect 9322 2986 9398 2996
rect 9034 2764 9110 2774
rect 9034 2708 9044 2764
rect 9100 2708 9110 2764
rect 9034 2698 9110 2708
rect 7594 2332 7670 2342
rect 7594 2276 7604 2332
rect 7660 2276 7670 2332
rect 7594 2266 7670 2276
rect 8890 2332 8966 2342
rect 8890 2276 8900 2332
rect 8956 2276 8966 2332
rect 8890 2266 8966 2276
rect 9042 2198 9102 2698
rect 9330 2486 9390 2986
rect 9322 2476 9398 2486
rect 9322 2420 9332 2476
rect 9388 2420 9398 2476
rect 9322 2410 9398 2420
rect 9474 2198 9534 3274
rect 9618 2342 9678 3706
rect 12930 3638 12990 3774
rect 13930 3772 14006 3782
rect 13930 3716 13940 3772
rect 13996 3716 14006 3772
rect 13930 3706 14006 3716
rect 14650 3772 14726 3782
rect 14650 3716 14660 3772
rect 14716 3716 14726 3772
rect 14650 3706 14726 3716
rect 10330 3628 10406 3638
rect 10330 3572 10340 3628
rect 10396 3572 10406 3628
rect 10330 3562 10406 3572
rect 10906 3628 10982 3638
rect 10906 3572 10916 3628
rect 10972 3572 10982 3628
rect 10906 3562 10982 3572
rect 12922 3628 12998 3638
rect 12922 3572 12932 3628
rect 12988 3572 12998 3628
rect 12922 3562 12998 3572
rect 13498 3628 13574 3638
rect 13498 3572 13508 3628
rect 13564 3572 13574 3628
rect 13498 3562 13574 3572
rect 9762 2774 9822 3342
rect 10186 3340 10262 3350
rect 10186 3284 10196 3340
rect 10252 3284 10262 3340
rect 10186 3274 10262 3284
rect 10194 2774 10254 3274
rect 10338 2918 10398 3562
rect 10762 3344 10838 3350
rect 10762 3280 10768 3344
rect 10832 3280 10838 3344
rect 10762 3274 10838 3280
rect 10330 2912 10406 2918
rect 10330 2848 10336 2912
rect 10400 2848 10406 2912
rect 10330 2842 10406 2848
rect 9754 2764 9830 2774
rect 9754 2708 9764 2764
rect 9820 2708 9830 2764
rect 9754 2698 9830 2708
rect 10186 2764 10262 2774
rect 10186 2708 10196 2764
rect 10252 2708 10262 2764
rect 10186 2698 10262 2708
rect 9762 2630 9822 2698
rect 9754 2620 9830 2630
rect 9754 2564 9764 2620
rect 9820 2564 9830 2620
rect 9754 2554 9830 2564
rect 10194 2342 10254 2698
rect 10338 2486 10398 2842
rect 10770 2774 10830 3274
rect 10914 3206 10974 3562
rect 12930 3350 12990 3562
rect 12058 3340 12134 3350
rect 12058 3284 12068 3340
rect 12124 3284 12134 3340
rect 12058 3274 12134 3284
rect 12922 3340 12998 3350
rect 12922 3284 12932 3340
rect 12988 3284 12998 3340
rect 12922 3274 12998 3284
rect 13210 3344 13286 3350
rect 13210 3280 13216 3344
rect 13280 3280 13286 3344
rect 13210 3274 13286 3280
rect 10906 3200 10982 3206
rect 10906 3136 10912 3200
rect 10976 3136 10982 3200
rect 10906 3130 10982 3136
rect 10762 2764 10838 2774
rect 10762 2708 10772 2764
rect 10828 2708 10838 2764
rect 10762 2698 10838 2708
rect 10914 2486 10974 3130
rect 12066 2774 12126 3274
rect 13218 2774 13278 3274
rect 13506 3206 13566 3562
rect 13498 3200 13574 3206
rect 13498 3136 13504 3200
rect 13568 3136 13574 3200
rect 13498 3130 13574 3136
rect 13506 2774 13566 3130
rect 11770 2768 11846 2774
rect 11770 2704 11776 2768
rect 11840 2704 11846 2768
rect 11770 2698 11846 2704
rect 12058 2764 12134 2774
rect 12058 2708 12068 2764
rect 12124 2708 12134 2764
rect 12058 2698 12134 2708
rect 13210 2764 13286 2774
rect 13210 2708 13220 2764
rect 13276 2708 13286 2764
rect 13210 2698 13286 2708
rect 13498 2764 13574 2774
rect 13498 2708 13508 2764
rect 13564 2708 13574 2764
rect 13498 2698 13574 2708
rect 10330 2476 10406 2486
rect 10330 2420 10340 2476
rect 10396 2420 10406 2476
rect 10330 2410 10406 2420
rect 10906 2476 10982 2486
rect 10906 2420 10916 2476
rect 10972 2420 10982 2476
rect 10906 2410 10982 2420
rect 9610 2332 9686 2342
rect 9610 2276 9620 2332
rect 9676 2276 9686 2332
rect 9610 2266 9686 2276
rect 10186 2332 10262 2342
rect 10186 2276 10196 2332
rect 10252 2276 10262 2332
rect 10186 2266 10262 2276
rect 4858 2188 4934 2198
rect 4858 2132 4868 2188
rect 4924 2132 4934 2188
rect 4858 2122 4934 2132
rect 5866 2188 5942 2198
rect 5866 2132 5876 2188
rect 5932 2132 5942 2188
rect 5866 2122 5942 2132
rect 6874 2188 6950 2198
rect 6874 2132 6884 2188
rect 6940 2132 6950 2188
rect 6874 2122 6950 2132
rect 9034 2188 9110 2198
rect 9034 2132 9044 2188
rect 9100 2132 9110 2188
rect 9034 2122 9110 2132
rect 9466 2188 9542 2198
rect 9466 2132 9476 2188
rect 9532 2132 9542 2188
rect 9466 2122 9542 2132
rect 2698 1904 2774 1910
rect 2698 1840 2704 1904
rect 2768 1840 2774 1904
rect 2698 1834 2774 1840
rect 5866 1904 5942 1910
rect 5866 1840 5872 1904
rect 5936 1840 5942 1904
rect 5866 1834 5942 1840
rect 6586 1900 6662 1910
rect 6586 1844 6596 1900
rect 6652 1844 6662 1900
rect 6586 1834 6662 1844
rect 7594 1900 7670 1910
rect 7594 1844 7604 1900
rect 7660 1844 7670 1900
rect 7594 1834 7670 1844
rect 8602 1900 8678 1910
rect 8602 1844 8612 1900
rect 8668 1844 8678 1900
rect 8602 1834 8678 1844
rect 10762 1900 10838 1910
rect 10762 1844 10772 1900
rect 10828 1844 10838 1900
rect 10762 1834 10838 1844
rect 11194 1900 11270 1910
rect 11194 1844 11204 1900
rect 11260 1844 11270 1900
rect 11194 1834 11270 1844
rect 3274 1756 3350 1766
rect 3274 1700 3284 1756
rect 3340 1700 3350 1756
rect 3274 1690 3350 1700
rect 826 1612 902 1622
rect 826 1556 836 1612
rect 892 1556 902 1612
rect 826 1546 902 1556
rect 682 1328 758 1334
rect 682 1264 688 1328
rect 752 1264 758 1328
rect 682 1258 758 1264
rect 690 758 750 1258
rect 834 1046 894 1546
rect 1402 1324 1478 1334
rect 1402 1268 1412 1324
rect 1468 1268 1478 1324
rect 1402 1258 1478 1268
rect 2554 1324 2630 1334
rect 2554 1268 2564 1324
rect 2620 1268 2630 1324
rect 2554 1258 2630 1268
rect 2842 1328 2918 1334
rect 2842 1264 2848 1328
rect 2912 1264 2918 1328
rect 2842 1258 2918 1264
rect 826 1036 902 1046
rect 826 980 836 1036
rect 892 980 902 1036
rect 826 970 902 980
rect 682 748 758 758
rect 682 692 692 748
rect 748 692 758 748
rect 682 682 758 692
rect 834 470 894 970
rect 1410 758 1470 1258
rect 2562 1046 2622 1258
rect 2554 1036 2630 1046
rect 2554 980 2564 1036
rect 2620 980 2630 1036
rect 2554 970 2630 980
rect 2562 758 2622 970
rect 1402 748 1478 758
rect 1402 692 1412 748
rect 1468 692 1478 748
rect 1402 682 1478 692
rect 2266 748 2342 758
rect 2266 692 2276 748
rect 2332 692 2342 748
rect 2266 682 2342 692
rect 2554 748 2630 758
rect 2554 692 2564 748
rect 2620 692 2630 748
rect 2554 682 2630 692
rect 2274 470 2334 682
rect 2850 470 2910 1258
rect 826 460 902 470
rect 826 404 836 460
rect 892 404 902 460
rect 826 394 902 404
rect 2266 460 2342 470
rect 2266 404 2276 460
rect 2332 404 2342 460
rect 2266 394 2342 404
rect 2842 460 2918 470
rect 2842 404 2852 460
rect 2908 404 2918 460
rect 2842 394 2918 404
rect 2274 258 2334 394
rect 3282 326 3342 1690
rect 4282 1612 4358 1622
rect 4282 1556 4292 1612
rect 4348 1556 4358 1612
rect 4282 1546 4358 1556
rect 4290 1334 4350 1546
rect 5874 1334 5934 1834
rect 6594 1622 6654 1834
rect 6010 1612 6086 1622
rect 6010 1556 6020 1612
rect 6076 1556 6086 1612
rect 6010 1546 6086 1556
rect 6586 1612 6662 1622
rect 6586 1556 6596 1612
rect 6652 1556 6662 1612
rect 6586 1546 6662 1556
rect 6018 1478 6078 1546
rect 6010 1468 6086 1478
rect 6010 1412 6020 1468
rect 6076 1412 6086 1468
rect 6010 1402 6086 1412
rect 6442 1468 6518 1478
rect 6442 1412 6452 1468
rect 6508 1412 6518 1468
rect 6442 1402 6518 1412
rect 3706 1324 3782 1334
rect 3706 1268 3716 1324
rect 3772 1268 3782 1324
rect 3706 1258 3782 1268
rect 3994 1324 4070 1334
rect 3994 1268 4004 1324
rect 4060 1268 4070 1324
rect 3994 1258 4070 1268
rect 4282 1328 4358 1334
rect 4282 1264 4288 1328
rect 4352 1264 4358 1328
rect 4282 1258 4358 1264
rect 5866 1324 5942 1334
rect 5866 1268 5876 1324
rect 5932 1268 5942 1324
rect 5866 1258 5942 1268
rect 3714 758 3774 1258
rect 4002 758 4062 1258
rect 3706 748 3782 758
rect 3706 692 3716 748
rect 3772 692 3782 748
rect 3706 682 3782 692
rect 3994 748 4070 758
rect 3994 692 4004 748
rect 4060 692 4070 748
rect 3994 682 4070 692
rect 4002 326 4062 682
rect 4290 470 4350 1258
rect 5874 758 5934 1258
rect 5866 748 5942 758
rect 5866 692 5876 748
rect 5932 692 5942 748
rect 5866 682 5942 692
rect 6018 470 6078 1402
rect 6450 1334 6510 1402
rect 6442 1324 6518 1334
rect 6442 1268 6452 1324
rect 6508 1268 6518 1324
rect 6442 1258 6518 1268
rect 6450 758 6510 1258
rect 6442 748 6518 758
rect 6442 692 6452 748
rect 6508 692 6518 748
rect 6442 682 6518 692
rect 6594 470 6654 1546
rect 7162 1328 7238 1334
rect 7162 1264 7168 1328
rect 7232 1264 7238 1328
rect 7162 1258 7238 1264
rect 7170 758 7230 1258
rect 7602 758 7662 1834
rect 7738 1756 7814 1766
rect 7738 1700 7748 1756
rect 7804 1700 7814 1756
rect 7738 1690 7814 1700
rect 8458 1756 8534 1766
rect 8458 1700 8468 1756
rect 8524 1700 8534 1756
rect 8458 1690 8534 1700
rect 7162 748 7238 758
rect 7162 692 7172 748
rect 7228 692 7238 748
rect 7162 682 7238 692
rect 7594 748 7670 758
rect 7594 692 7604 748
rect 7660 692 7670 748
rect 7594 682 7670 692
rect 4282 460 4358 470
rect 4282 404 4292 460
rect 4348 404 4358 460
rect 4282 394 4358 404
rect 6010 460 6086 470
rect 6010 404 6020 460
rect 6076 404 6086 460
rect 6010 394 6086 404
rect 6586 460 6662 470
rect 6586 404 6596 460
rect 6652 404 6662 460
rect 6586 394 6662 404
rect 7746 326 7806 1690
rect 7882 1468 7958 1478
rect 7882 1412 7892 1468
rect 7948 1412 7958 1468
rect 7882 1402 7958 1412
rect 8314 1468 8390 1478
rect 8314 1412 8324 1468
rect 8380 1412 8390 1468
rect 8314 1402 8390 1412
rect 7890 1334 7950 1402
rect 7882 1324 7958 1334
rect 7882 1268 7892 1324
rect 7948 1268 7958 1324
rect 7882 1258 7958 1268
rect 7890 690 7950 1258
rect 8178 1046 8238 1326
rect 8170 1036 8246 1046
rect 8170 980 8180 1036
rect 8236 980 8246 1036
rect 8170 970 8246 980
rect 8178 690 8238 970
rect 8322 758 8382 1402
rect 8314 748 8390 758
rect 8314 692 8324 748
rect 8380 692 8390 748
rect 8314 682 8390 692
rect 8466 326 8526 1690
rect 8610 1334 8670 1834
rect 9322 1756 9398 1766
rect 9322 1700 9332 1756
rect 9388 1700 9398 1756
rect 9322 1690 9398 1700
rect 10618 1756 10694 1766
rect 10618 1700 10628 1756
rect 10684 1700 10694 1756
rect 10618 1690 10694 1700
rect 9330 1334 9390 1690
rect 9466 1612 9542 1622
rect 9466 1556 9476 1612
rect 9532 1556 9542 1612
rect 9466 1546 9542 1556
rect 8602 1324 8678 1334
rect 8602 1268 8612 1324
rect 8668 1268 8678 1324
rect 8602 1258 8678 1268
rect 9322 1324 9398 1334
rect 9322 1268 9332 1324
rect 9388 1268 9398 1324
rect 9322 1258 9398 1268
rect 8610 690 8670 1258
rect 9330 758 9390 1258
rect 9474 1046 9534 1546
rect 10474 1468 10550 1478
rect 10474 1412 10484 1468
rect 10540 1412 10550 1468
rect 10474 1402 10550 1412
rect 10042 1324 10118 1334
rect 10042 1268 10052 1324
rect 10108 1268 10118 1324
rect 10042 1258 10118 1268
rect 10050 1046 10110 1258
rect 9466 1036 9542 1046
rect 9466 980 9476 1036
rect 9532 980 9542 1036
rect 9466 970 9542 980
rect 10042 1036 10118 1046
rect 10042 980 10052 1036
rect 10108 980 10118 1036
rect 10042 970 10118 980
rect 9322 748 9398 758
rect 9322 692 9332 748
rect 9388 692 9398 748
rect 9322 682 9398 692
rect 9474 470 9534 970
rect 10050 758 10110 970
rect 10482 758 10542 1402
rect 10042 748 10118 758
rect 10042 692 10052 748
rect 10108 692 10118 748
rect 10042 682 10118 692
rect 10474 748 10550 758
rect 10474 692 10484 748
rect 10540 692 10550 748
rect 10474 682 10550 692
rect 9466 460 9542 470
rect 9466 404 9476 460
rect 9532 404 9542 460
rect 9466 394 9542 404
rect 10626 326 10686 1690
rect 10770 1334 10830 1834
rect 11050 1612 11126 1622
rect 11050 1556 11060 1612
rect 11116 1556 11126 1612
rect 11050 1546 11126 1556
rect 10762 1324 10838 1334
rect 10762 1268 10772 1324
rect 10828 1268 10838 1324
rect 10762 1258 10838 1268
rect 10770 690 10830 1258
rect 11058 1046 11118 1546
rect 11050 1036 11126 1046
rect 11050 980 11060 1036
rect 11116 980 11126 1036
rect 11050 970 11126 980
rect 11058 690 11118 970
rect 11202 758 11262 1834
rect 11338 1756 11414 1766
rect 11338 1700 11348 1756
rect 11404 1700 11414 1756
rect 11338 1690 11414 1700
rect 11194 748 11270 758
rect 11194 692 11204 748
rect 11260 692 11270 748
rect 11194 682 11270 692
rect 11346 326 11406 1690
rect 11482 1468 11558 1478
rect 11482 1412 11492 1468
rect 11548 1412 11558 1468
rect 11482 1402 11558 1412
rect 11490 1334 11550 1402
rect 11778 1334 11838 2698
rect 13938 2342 13998 3706
rect 14658 3350 14718 3706
rect 14938 3628 15014 3638
rect 14938 3572 14948 3628
rect 15004 3572 15014 3628
rect 14938 3562 15014 3572
rect 16666 3628 16742 3638
rect 16666 3572 16676 3628
rect 16732 3572 16742 3628
rect 16666 3562 16742 3572
rect 14362 3340 14438 3350
rect 14362 3284 14372 3340
rect 14428 3284 14438 3340
rect 14362 3274 14438 3284
rect 14650 3340 14726 3350
rect 14650 3284 14660 3340
rect 14716 3284 14726 3340
rect 14650 3274 14726 3284
rect 14370 2918 14430 3274
rect 14362 2912 14438 2918
rect 14362 2848 14368 2912
rect 14432 2848 14438 2912
rect 14362 2842 14438 2848
rect 14370 2774 14430 2842
rect 14658 2774 14718 3274
rect 14362 2764 14438 2774
rect 14362 2708 14372 2764
rect 14428 2708 14438 2764
rect 14362 2698 14438 2708
rect 14650 2764 14726 2774
rect 14650 2708 14660 2764
rect 14716 2708 14726 2764
rect 14650 2698 14726 2708
rect 14946 2486 15006 3562
rect 16674 2486 16734 3562
rect 19978 3340 20054 3350
rect 19978 3284 19988 3340
rect 20044 3284 20054 3340
rect 19978 3274 20054 3284
rect 19986 2774 20046 3274
rect 19978 2764 20054 2774
rect 19978 2708 19988 2764
rect 20044 2708 20054 2764
rect 19978 2698 20054 2708
rect 19986 2630 20046 2698
rect 19978 2624 20054 2630
rect 19978 2560 19984 2624
rect 20048 2560 20054 2624
rect 19978 2554 20054 2560
rect 20698 2624 20774 2630
rect 20698 2560 20704 2624
rect 20768 2560 20774 2624
rect 20698 2554 20774 2560
rect 14938 2476 15014 2486
rect 14938 2420 14948 2476
rect 15004 2420 15014 2476
rect 14938 2410 15014 2420
rect 16666 2476 16742 2486
rect 16666 2420 16676 2476
rect 16732 2420 16742 2476
rect 16666 2410 16742 2420
rect 13930 2332 14006 2342
rect 13930 2276 13940 2332
rect 13996 2276 14006 2332
rect 13930 2266 14006 2276
rect 14946 2198 15006 2410
rect 14650 2192 14726 2198
rect 14650 2128 14656 2192
rect 14720 2128 14726 2192
rect 14650 2122 14726 2128
rect 14938 2192 15014 2198
rect 14938 2128 14944 2192
rect 15008 2128 15014 2192
rect 14938 2122 15014 2128
rect 11914 1756 11990 1766
rect 11914 1700 11924 1756
rect 11980 1700 11990 1756
rect 11914 1690 11990 1700
rect 11922 1334 11982 1690
rect 12058 1612 12134 1622
rect 12058 1556 12068 1612
rect 12124 1556 12134 1612
rect 12058 1546 12134 1556
rect 12634 1612 12710 1622
rect 12634 1556 12644 1612
rect 12700 1556 12710 1612
rect 12634 1546 12710 1556
rect 13210 1612 13286 1622
rect 13210 1556 13220 1612
rect 13276 1556 13286 1612
rect 13210 1546 13286 1556
rect 13786 1612 13862 1622
rect 13786 1556 13796 1612
rect 13852 1556 13862 1612
rect 13786 1546 13862 1556
rect 12066 1334 12126 1546
rect 11482 1324 11558 1334
rect 11482 1268 11492 1324
rect 11548 1268 11558 1324
rect 11482 1258 11558 1268
rect 11770 1328 11846 1334
rect 11770 1264 11776 1328
rect 11840 1264 11846 1328
rect 11770 1258 11846 1264
rect 11914 1324 11990 1334
rect 11914 1268 11924 1324
rect 11980 1268 11990 1324
rect 11914 1258 11990 1268
rect 12058 1328 12134 1334
rect 12058 1264 12064 1328
rect 12128 1264 12134 1328
rect 12058 1258 12134 1264
rect 12490 1328 12566 1334
rect 12490 1264 12496 1328
rect 12560 1264 12566 1328
rect 12490 1258 12566 1264
rect 11490 690 11550 1258
rect 11922 758 11982 1258
rect 11914 748 11990 758
rect 11914 692 11924 748
rect 11980 692 11990 748
rect 11914 682 11990 692
rect 12066 470 12126 1258
rect 12498 758 12558 1258
rect 12642 1046 12702 1546
rect 13218 1334 13278 1546
rect 13066 1324 13142 1334
rect 13066 1268 13076 1324
rect 13132 1268 13142 1324
rect 13066 1258 13142 1268
rect 13210 1328 13286 1334
rect 13210 1264 13216 1328
rect 13280 1264 13286 1328
rect 13210 1258 13286 1264
rect 13642 1328 13718 1334
rect 13642 1264 13648 1328
rect 13712 1264 13718 1328
rect 13642 1258 13718 1264
rect 13074 1046 13134 1258
rect 12634 1036 12710 1046
rect 12634 980 12644 1036
rect 12700 980 12710 1036
rect 12634 970 12710 980
rect 13066 1036 13142 1046
rect 13066 980 13076 1036
rect 13132 980 13142 1036
rect 13066 970 13142 980
rect 12490 748 12566 758
rect 12490 692 12500 748
rect 12556 692 12566 748
rect 12490 682 12566 692
rect 12642 470 12702 970
rect 13074 758 13134 970
rect 13066 748 13142 758
rect 13066 692 13076 748
rect 13132 692 13142 748
rect 13066 682 13142 692
rect 13218 470 13278 1258
rect 13650 758 13710 1258
rect 13794 1046 13854 1546
rect 14658 1334 14718 2122
rect 20706 1622 20766 2554
rect 14938 1612 15014 1622
rect 14938 1556 14948 1612
rect 15004 1556 15014 1612
rect 14938 1546 15014 1556
rect 15514 1612 15590 1622
rect 15514 1556 15524 1612
rect 15580 1556 15590 1612
rect 15514 1546 15590 1556
rect 16378 1612 16454 1622
rect 16378 1556 16388 1612
rect 16444 1556 16454 1612
rect 16378 1546 16454 1556
rect 20698 1612 20774 1622
rect 20698 1556 20708 1612
rect 20764 1556 20774 1612
rect 20698 1546 20774 1556
rect 14650 1328 14726 1334
rect 14650 1264 14656 1328
rect 14720 1264 14726 1328
rect 14650 1258 14726 1264
rect 14794 1324 14870 1334
rect 14794 1268 14804 1324
rect 14860 1268 14870 1324
rect 14794 1258 14870 1268
rect 14802 1046 14862 1258
rect 13786 1036 13862 1046
rect 13786 980 13796 1036
rect 13852 980 13862 1036
rect 13786 970 13862 980
rect 14794 1036 14870 1046
rect 14794 980 14804 1036
rect 14860 980 14870 1036
rect 14794 970 14870 980
rect 13642 748 13718 758
rect 13642 692 13652 748
rect 13708 692 13718 748
rect 13642 682 13718 692
rect 13794 470 13854 970
rect 14802 758 14862 970
rect 14794 748 14870 758
rect 14794 692 14804 748
rect 14860 692 14870 748
rect 14794 682 14870 692
rect 14946 470 15006 1546
rect 15522 1190 15582 1546
rect 16386 1334 16446 1546
rect 15658 1328 15734 1334
rect 15658 1264 15664 1328
rect 15728 1264 15734 1328
rect 15658 1258 15734 1264
rect 15946 1324 16022 1334
rect 15946 1268 15956 1324
rect 16012 1268 16022 1324
rect 15946 1258 16022 1268
rect 16378 1328 16454 1334
rect 16378 1264 16384 1328
rect 16448 1264 16454 1328
rect 16378 1258 16454 1264
rect 17386 1328 17462 1334
rect 17386 1264 17392 1328
rect 17456 1264 17462 1328
rect 17386 1258 17462 1264
rect 15514 1184 15590 1190
rect 15514 1120 15520 1184
rect 15584 1120 15590 1184
rect 15514 1114 15590 1120
rect 15522 470 15582 1114
rect 15666 758 15726 1258
rect 15954 1190 16014 1258
rect 15946 1184 16022 1190
rect 15946 1120 15952 1184
rect 16016 1120 16022 1184
rect 15946 1114 16022 1120
rect 15954 758 16014 1114
rect 15658 748 15734 758
rect 15658 692 15668 748
rect 15724 692 15734 748
rect 15658 682 15734 692
rect 15946 748 16022 758
rect 15946 692 15956 748
rect 16012 692 16022 748
rect 15946 682 16022 692
rect 16386 470 16446 1258
rect 17394 758 17454 1258
rect 17386 748 17462 758
rect 17386 692 17396 748
rect 17452 692 17462 748
rect 17386 682 17462 692
rect 20706 470 20766 1546
rect 12058 460 12134 470
rect 12058 404 12068 460
rect 12124 404 12134 460
rect 12058 394 12134 404
rect 12634 460 12710 470
rect 12634 404 12644 460
rect 12700 404 12710 460
rect 12634 394 12710 404
rect 13210 460 13286 470
rect 13210 404 13220 460
rect 13276 404 13286 460
rect 13210 394 13286 404
rect 13786 460 13862 470
rect 13786 404 13796 460
rect 13852 404 13862 460
rect 13786 394 13862 404
rect 14938 460 15014 470
rect 14938 404 14948 460
rect 15004 404 15014 460
rect 14938 394 15014 404
rect 15514 460 15590 470
rect 15514 404 15524 460
rect 15580 404 15590 460
rect 15514 394 15590 404
rect 16378 460 16454 470
rect 16378 404 16388 460
rect 16444 404 16454 460
rect 16378 394 16454 404
rect 20698 460 20774 470
rect 20698 404 20708 460
rect 20764 404 20774 460
rect 20698 394 20774 404
rect 3274 316 3350 326
rect 3274 260 3284 316
rect 3340 260 3350 316
rect 3274 250 3350 260
rect 3994 316 4070 326
rect 3994 260 4004 316
rect 4060 260 4070 316
rect 3994 250 4070 260
rect 7738 316 7814 326
rect 7738 260 7748 316
rect 7804 260 7814 316
rect 7738 250 7814 260
rect 8458 316 8534 326
rect 8458 260 8468 316
rect 8524 260 8534 316
rect 8458 250 8534 260
rect 10618 316 10694 326
rect 10618 260 10628 316
rect 10684 260 10694 316
rect 10618 250 10694 260
rect 11338 316 11414 326
rect 11338 260 11348 316
rect 11404 260 11414 316
rect 11338 250 11414 260
<< via3 >>
rect 976 2764 1040 2768
rect 976 2708 980 2764
rect 980 2708 1036 2764
rect 1036 2708 1040 2764
rect 976 2704 1040 2708
rect 1408 2704 1472 2768
rect 2128 2764 2192 2768
rect 2128 2708 2132 2764
rect 2132 2708 2188 2764
rect 2188 2708 2192 2764
rect 2128 2704 2192 2708
rect 2560 2704 2624 2768
rect 3136 2704 3200 2768
rect 4144 2764 4208 2768
rect 4144 2708 4148 2764
rect 4148 2708 4204 2764
rect 4204 2708 4208 2764
rect 4144 2704 4208 2708
rect 5440 2764 5504 2768
rect 5440 2708 5444 2764
rect 5444 2708 5500 2764
rect 5500 2708 5504 2764
rect 5440 2704 5504 2708
rect 10768 3340 10832 3344
rect 10768 3284 10772 3340
rect 10772 3284 10828 3340
rect 10828 3284 10832 3340
rect 10768 3280 10832 3284
rect 10336 2848 10400 2912
rect 13216 3340 13280 3344
rect 13216 3284 13220 3340
rect 13220 3284 13276 3340
rect 13276 3284 13280 3340
rect 13216 3280 13280 3284
rect 10912 3136 10976 3200
rect 13504 3136 13568 3200
rect 11776 2704 11840 2768
rect 2704 1840 2768 1904
rect 5872 1840 5936 1904
rect 688 1324 752 1328
rect 688 1268 692 1324
rect 692 1268 748 1324
rect 748 1268 752 1324
rect 688 1264 752 1268
rect 2848 1324 2912 1328
rect 2848 1268 2852 1324
rect 2852 1268 2908 1324
rect 2908 1268 2912 1324
rect 2848 1264 2912 1268
rect 4288 1264 4352 1328
rect 7168 1324 7232 1328
rect 7168 1268 7172 1324
rect 7172 1268 7228 1324
rect 7228 1268 7232 1324
rect 7168 1264 7232 1268
rect 14368 2848 14432 2912
rect 19984 2560 20048 2624
rect 20704 2560 20768 2624
rect 14656 2128 14720 2192
rect 14944 2128 15008 2192
rect 11776 1264 11840 1328
rect 12064 1264 12128 1328
rect 12496 1324 12560 1328
rect 12496 1268 12500 1324
rect 12500 1268 12556 1324
rect 12556 1268 12560 1324
rect 12496 1264 12560 1268
rect 13216 1264 13280 1328
rect 13648 1324 13712 1328
rect 13648 1268 13652 1324
rect 13652 1268 13708 1324
rect 13708 1268 13712 1324
rect 13648 1264 13712 1268
rect 14656 1264 14720 1328
rect 15664 1324 15728 1328
rect 15664 1268 15668 1324
rect 15668 1268 15724 1324
rect 15724 1268 15728 1324
rect 15664 1264 15728 1268
rect 16384 1264 16448 1328
rect 17392 1324 17456 1328
rect 17392 1268 17396 1324
rect 17396 1268 17452 1324
rect 17452 1268 17456 1324
rect 17392 1264 17456 1268
rect 15520 1120 15584 1184
rect 15952 1120 16016 1184
<< metal4 >>
rect 10766 3344 10834 3346
rect 10766 3280 10768 3344
rect 10832 3342 10834 3344
rect 13214 3344 13282 3346
rect 13214 3342 13216 3344
rect 10832 3282 13216 3342
rect 10832 3280 10834 3282
rect 10766 3278 10834 3280
rect 13214 3280 13216 3282
rect 13280 3280 13282 3344
rect 13214 3278 13282 3280
rect 10910 3200 10978 3202
rect 10910 3136 10912 3200
rect 10976 3198 10978 3200
rect 13502 3200 13570 3202
rect 13502 3198 13504 3200
rect 10976 3138 13504 3198
rect 10976 3136 10978 3138
rect 10910 3134 10978 3136
rect 13502 3136 13504 3138
rect 13568 3136 13570 3200
rect 13502 3134 13570 3136
rect 10334 2912 10402 2914
rect 10334 2848 10336 2912
rect 10400 2910 10402 2912
rect 14366 2912 14434 2914
rect 14366 2910 14368 2912
rect 10400 2850 14368 2910
rect 10400 2848 10402 2850
rect 10334 2846 10402 2848
rect 14366 2848 14368 2850
rect 14432 2848 14434 2912
rect 14366 2846 14434 2848
rect 974 2768 1042 2770
rect 974 2704 976 2768
rect 1040 2766 1042 2768
rect 1406 2768 1474 2770
rect 1406 2766 1408 2768
rect 1040 2706 1408 2766
rect 1040 2704 1042 2706
rect 974 2702 1042 2704
rect 1406 2704 1408 2706
rect 1472 2704 1474 2768
rect 1406 2702 1474 2704
rect 2126 2768 2194 2770
rect 2126 2704 2128 2768
rect 2192 2766 2194 2768
rect 2558 2768 2626 2770
rect 2558 2766 2560 2768
rect 2192 2706 2560 2766
rect 2192 2704 2194 2706
rect 2126 2702 2194 2704
rect 2558 2704 2560 2706
rect 2624 2704 2626 2768
rect 2558 2702 2626 2704
rect 3134 2768 3202 2770
rect 3134 2704 3136 2768
rect 3200 2766 3202 2768
rect 4142 2768 4210 2770
rect 4142 2766 4144 2768
rect 3200 2706 4144 2766
rect 3200 2704 3202 2706
rect 3134 2702 3202 2704
rect 4142 2704 4144 2706
rect 4208 2704 4210 2768
rect 4142 2702 4210 2704
rect 5438 2768 5506 2770
rect 5438 2704 5440 2768
rect 5504 2766 5506 2768
rect 11774 2768 11842 2770
rect 11774 2766 11776 2768
rect 5504 2706 11776 2766
rect 5504 2704 5506 2706
rect 5438 2702 5506 2704
rect 11774 2704 11776 2706
rect 11840 2704 11842 2768
rect 11774 2702 11842 2704
rect 19982 2624 20050 2626
rect 19982 2560 19984 2624
rect 20048 2622 20050 2624
rect 20702 2624 20770 2626
rect 20702 2622 20704 2624
rect 20048 2562 20704 2622
rect 20048 2560 20050 2562
rect 19982 2558 20050 2560
rect 20702 2560 20704 2562
rect 20768 2560 20770 2624
rect 20702 2558 20770 2560
rect 14654 2192 14722 2194
rect 14654 2128 14656 2192
rect 14720 2190 14722 2192
rect 14942 2192 15010 2194
rect 14942 2190 14944 2192
rect 14720 2130 14944 2190
rect 14720 2128 14722 2130
rect 14654 2126 14722 2128
rect 14942 2128 14944 2130
rect 15008 2128 15010 2192
rect 14942 2126 15010 2128
rect 2702 1904 2770 1906
rect 2702 1840 2704 1904
rect 2768 1902 2770 1904
rect 5870 1904 5938 1906
rect 5870 1902 5872 1904
rect 2768 1842 5872 1902
rect 2768 1840 2770 1842
rect 2702 1838 2770 1840
rect 5870 1840 5872 1842
rect 5936 1840 5938 1904
rect 5870 1838 5938 1840
rect 686 1328 754 1330
rect 686 1264 688 1328
rect 752 1326 754 1328
rect 2846 1328 2914 1330
rect 2846 1326 2848 1328
rect 752 1266 2848 1326
rect 752 1264 754 1266
rect 686 1262 754 1264
rect 2846 1264 2848 1266
rect 2912 1264 2914 1328
rect 2846 1262 2914 1264
rect 4286 1328 4354 1330
rect 4286 1264 4288 1328
rect 4352 1326 4354 1328
rect 7166 1328 7234 1330
rect 7166 1326 7168 1328
rect 4352 1266 7168 1326
rect 4352 1264 4354 1266
rect 4286 1262 4354 1264
rect 7166 1264 7168 1266
rect 7232 1264 7234 1328
rect 7166 1262 7234 1264
rect 11774 1328 11842 1330
rect 11774 1264 11776 1328
rect 11840 1326 11842 1328
rect 12062 1328 12130 1330
rect 12062 1326 12064 1328
rect 11840 1266 12064 1326
rect 11840 1264 11842 1266
rect 11774 1262 11842 1264
rect 12062 1264 12064 1266
rect 12128 1326 12130 1328
rect 12494 1328 12562 1330
rect 12494 1326 12496 1328
rect 12128 1266 12496 1326
rect 12128 1264 12130 1266
rect 12062 1262 12130 1264
rect 12494 1264 12496 1266
rect 12560 1264 12562 1328
rect 12494 1262 12562 1264
rect 13214 1328 13282 1330
rect 13214 1264 13216 1328
rect 13280 1326 13282 1328
rect 13646 1328 13714 1330
rect 13646 1326 13648 1328
rect 13280 1266 13648 1326
rect 13280 1264 13282 1266
rect 13214 1262 13282 1264
rect 13646 1264 13648 1266
rect 13712 1264 13714 1328
rect 13646 1262 13714 1264
rect 14654 1328 14722 1330
rect 14654 1264 14656 1328
rect 14720 1326 14722 1328
rect 15662 1328 15730 1330
rect 15662 1326 15664 1328
rect 14720 1266 15664 1326
rect 14720 1264 14722 1266
rect 14654 1262 14722 1264
rect 15662 1264 15664 1266
rect 15728 1264 15730 1328
rect 15662 1262 15730 1264
rect 16382 1328 16450 1330
rect 16382 1264 16384 1328
rect 16448 1326 16450 1328
rect 17390 1328 17458 1330
rect 17390 1326 17392 1328
rect 16448 1266 17392 1326
rect 16448 1264 16450 1266
rect 16382 1262 16450 1264
rect 17390 1264 17392 1266
rect 17456 1264 17458 1328
rect 17390 1262 17458 1264
rect 15518 1184 15586 1186
rect 15518 1120 15520 1184
rect 15584 1182 15586 1184
rect 15950 1184 16018 1186
rect 15950 1182 15952 1184
rect 15584 1122 15952 1182
rect 15584 1120 15586 1122
rect 15518 1118 15586 1120
rect 15950 1120 15952 1122
rect 16016 1120 16018 1184
rect 15950 1118 16018 1120
<< labels >>
flabel metal3 2736 3024 2736 3024 0 FreeSans 480 90 0 0 SCAN_CLK
port 1 nsew
flabel metal3 864 3024 864 3024 0 FreeSans 480 90 0 0 SCAN_CLK_OUT
port 2 nsew
flabel metal3 3744 1008 3744 1008 0 FreeSans 480 90 0 0 SCAN_DATA_IN
port 3 nsew
flabel metal3 16704 3024 16704 3024 0 FreeSans 480 90 0 0 SCAN_DATA_OUT
port 4 nsew
flabel metal3 3024 3024 3024 3024 0 FreeSans 480 90 0 0 SCAN_EN
port 5 nsew
flabel metal3 13248 3024 13248 3024 0 FreeSans 480 90 0 0 SCAN_GATE
port 6 nsew
flabel metal3 12096 3024 12096 3024 0 FreeSans 480 90 0 0 SCAN_GATE_VALUE
port 7 nsew
flabel metal3 1440 1008 1440 1008 0 FreeSans 480 90 0 0 SCAN_IN
port 8 nsew
flabel metal3 720 1008 720 1008 0 FreeSans 480 90 0 0 SCAN_LOAD
port 9 nsew
flabel metal3 14976 1008 14976 1008 0 FreeSans 480 90 0 0 SCAN_OUT
port 10 nsew
flabel metal2 10512 0 10512 0 0 FreeSans 960 0 0 0 VDD_
port 11 nsew
flabel metal2 10512 4032 10512 4032 0 FreeSans 960 0 0 0 VDD_
port 12 nsew
flabel metal2 10512 2016 10512 2016 0 FreeSans 960 0 0 0 VSS
port 13 nsew
flabel metal3 720 1008 720 1008 0 FreeSans 480 90 0 0 I0/I
flabel metal3 864 1008 864 1008 0 FreeSans 480 90 0 0 I0/O
flabel metal2 864 2016 864 2016 0 FreeSans 960 0 0 0 I0/VSS
flabel metal2 864 0 864 0 0 FreeSans 960 0 0 0 I0/VDD
flabel metal1 834 188 894 594 0 FreeSans 160 0 0 0 I0/MP0_IM0/D0
flabel metal1 776 684 950 756 0 FreeSans 160 0 0 0 I0/MP0_IM0/G0
flabel metal1 690 188 750 594 0 FreeSans 160 0 0 0 I0/MP0_IM0/S0
flabel metal1 978 188 1038 594 0 FreeSans 160 0 0 0 I0/MP0_IM0/S1
flabel nwell 700 654 724 670 0 FreeSans 80 0 0 0 I0/MP0_IM0/BODY
flabel space 1008 0 1152 1008 0 FreeSans 320 90 0 0 I0/MP0_IBNDR0/pmos_boundary
flabel space 576 0 720 1008 0 FreeSans 320 90 0 0 I0/MP0_IBNDL0/pmos_boundary
flabel metal1 690 1402 750 1728 0 FreeSans 240 0 0 0 I0/MN0_IM0/S0
flabel metal1 834 1402 894 1728 0 FreeSans 240 0 0 0 I0/MN0_IM0/D0
flabel metal1 978 1402 1038 1728 0 FreeSans 240 0 0 0 I0/MN0_IM0/S1
flabel metal1 776 1260 950 1332 0 FreeSans 240 0 0 0 I0/MN0_IM0/G0
rlabel pwell 680 1340 710 1362 5 I0/MN0_IM0/BODY
flabel space 1008 1008 1152 2016 0 FreeSans 320 90 0 0 I0/MN0_IBNDR0/nmos_boundary
flabel space 576 1008 720 2016 0 FreeSans 320 90 0 0 I0/MN0_IBNDL0/nmos_boundary
flabel metal3 1008 3024 1008 3024 0 FreeSans 480 90 0 0 I15/I
flabel metal3 864 3024 864 3024 0 FreeSans 480 90 0 0 I15/O
flabel metal2 864 2016 864 2016 0 FreeSans 960 0 0 0 I15/VSS
flabel metal2 864 4032 864 4032 0 FreeSans 960 0 0 0 I15/VDD
flabel metal1 834 3438 894 3844 0 FreeSans 160 0 0 0 I15/MP0_IM0/D0
flabel metal1 778 3276 952 3348 0 FreeSans 160 0 0 0 I15/MP0_IM0/G0
flabel metal1 978 3438 1038 3844 0 FreeSans 160 0 0 0 I15/MP0_IM0/S0
flabel metal1 690 3438 750 3844 0 FreeSans 160 0 0 0 I15/MP0_IM0/S1
flabel nwell 1004 3362 1028 3378 0 FreeSans 80 0 0 0 I15/MP0_IM0/BODY
flabel space 576 3024 720 4032 0 FreeSans 320 90 0 0 I15/MP0_IBNDR0/pmos_boundary
flabel space 1008 3024 1152 4032 0 FreeSans 320 90 0 0 I15/MP0_IBNDL0/pmos_boundary
flabel metal1 978 2304 1038 2630 0 FreeSans 240 0 0 0 I15/MN0_IM0/S0
flabel metal1 834 2304 894 2630 0 FreeSans 240 0 0 0 I15/MN0_IM0/D0
flabel metal1 690 2304 750 2630 0 FreeSans 240 0 0 0 I15/MN0_IM0/S1
flabel metal1 778 2700 952 2772 0 FreeSans 240 0 0 0 I15/MN0_IM0/G0
rlabel pwell 1018 2670 1048 2692 1 I15/MN0_IM0/BODY
flabel space 576 2016 720 3024 0 FreeSans 320 90 0 0 I15/MN0_IBNDR0/nmos_boundary
flabel space 1008 2016 1152 3024 0 FreeSans 320 90 0 0 I15/MN0_IBNDL0/nmos_boundary
flabel space 432 0 576 1024 0 FreeSans 320 90 0 0 TAP0_0/MPT0_IBNDR0/ptap_boundary
flabel space 0 0 144 1024 0 FreeSans 320 90 0 0 TAP0_0/MPT0_IBNDL0/ptap_boundary
flabel space 432 992 576 2016 0 FreeSans 320 90 0 0 TAP0_0/MNT0_IBNDR0/ntap_boundary
flabel space 0 992 144 2016 0 FreeSans 320 90 0 0 TAP0_0/MNT0_IBNDL0/ntap_boundary
flabel space 432 3008 576 4032 0 FreeSans 320 90 0 0 TAP1_0/MPT0_IBNDR0/ptap_boundary
flabel space 0 3008 144 4032 0 FreeSans 320 90 0 0 TAP1_0/MPT0_IBNDL0/ptap_boundary
flabel space 432 2016 576 3040 0 FreeSans 320 90 0 0 TAP1_0/MNT0_IBNDR0/ntap_boundary
flabel space 0 2016 144 3040 0 FreeSans 320 90 0 0 TAP1_0/MNT0_IBNDL0/ntap_boundary
flabel metal3 1584 3024 1584 3024 0 FreeSans 480 90 0 0 I16/I
flabel metal3 1440 3024 1440 3024 0 FreeSans 480 90 0 0 I16/O
flabel metal2 1440 2016 1440 2016 0 FreeSans 960 0 0 0 I16/VSS
flabel metal2 1440 4032 1440 4032 0 FreeSans 960 0 0 0 I16/VDD
flabel metal1 1410 3438 1470 3844 0 FreeSans 160 0 0 0 I16/MP0_IM0/D0
flabel metal1 1354 3276 1528 3348 0 FreeSans 160 0 0 0 I16/MP0_IM0/G0
flabel metal1 1554 3438 1614 3844 0 FreeSans 160 0 0 0 I16/MP0_IM0/S0
flabel metal1 1266 3438 1326 3844 0 FreeSans 160 0 0 0 I16/MP0_IM0/S1
flabel nwell 1580 3362 1604 3378 0 FreeSans 80 0 0 0 I16/MP0_IM0/BODY
flabel space 1152 3024 1296 4032 0 FreeSans 320 90 0 0 I16/MP0_IBNDR0/pmos_boundary
flabel space 1584 3024 1728 4032 0 FreeSans 320 90 0 0 I16/MP0_IBNDL0/pmos_boundary
flabel metal1 1554 2304 1614 2630 0 FreeSans 240 0 0 0 I16/MN0_IM0/S0
flabel metal1 1410 2304 1470 2630 0 FreeSans 240 0 0 0 I16/MN0_IM0/D0
flabel metal1 1266 2304 1326 2630 0 FreeSans 240 0 0 0 I16/MN0_IM0/S1
flabel metal1 1354 2700 1528 2772 0 FreeSans 240 0 0 0 I16/MN0_IM0/G0
rlabel pwell 1594 2670 1624 2692 1 I16/MN0_IM0/BODY
flabel space 1152 2016 1296 3024 0 FreeSans 320 90 0 0 I16/MN0_IBNDR0/nmos_boundary
flabel space 1584 2016 1728 3024 0 FreeSans 320 90 0 0 I16/MN0_IBNDL0/nmos_boundary
flabel metal3 2160 3024 2160 3024 0 FreeSans 480 90 0 0 I17/I
flabel metal3 2016 3024 2016 3024 0 FreeSans 480 90 0 0 I17/O
flabel metal2 2016 2016 2016 2016 0 FreeSans 960 0 0 0 I17/VSS
flabel metal2 2016 4032 2016 4032 0 FreeSans 960 0 0 0 I17/VDD
flabel metal1 1986 3438 2046 3844 0 FreeSans 160 0 0 0 I17/MP0_IM0/D0
flabel metal1 1930 3276 2104 3348 0 FreeSans 160 0 0 0 I17/MP0_IM0/G0
flabel metal1 2130 3438 2190 3844 0 FreeSans 160 0 0 0 I17/MP0_IM0/S0
flabel metal1 1842 3438 1902 3844 0 FreeSans 160 0 0 0 I17/MP0_IM0/S1
flabel nwell 2156 3362 2180 3378 0 FreeSans 80 0 0 0 I17/MP0_IM0/BODY
flabel space 1728 3024 1872 4032 0 FreeSans 320 90 0 0 I17/MP0_IBNDR0/pmos_boundary
flabel space 2160 3024 2304 4032 0 FreeSans 320 90 0 0 I17/MP0_IBNDL0/pmos_boundary
flabel metal1 2130 2304 2190 2630 0 FreeSans 240 0 0 0 I17/MN0_IM0/S0
flabel metal1 1986 2304 2046 2630 0 FreeSans 240 0 0 0 I17/MN0_IM0/D0
flabel metal1 1842 2304 1902 2630 0 FreeSans 240 0 0 0 I17/MN0_IM0/S1
flabel metal1 1930 2700 2104 2772 0 FreeSans 240 0 0 0 I17/MN0_IM0/G0
rlabel pwell 2170 2670 2200 2692 1 I17/MN0_IM0/BODY
flabel space 1728 2016 1872 3024 0 FreeSans 320 90 0 0 I17/MN0_IBNDR0/nmos_boundary
flabel space 2160 2016 2304 3024 0 FreeSans 320 90 0 0 I17/MN0_IBNDL0/nmos_boundary
flabel metal3 2736 3024 2736 3024 0 FreeSans 480 90 0 0 I18/I
flabel metal3 2592 3024 2592 3024 0 FreeSans 480 90 0 0 I18/O
flabel metal2 2592 2016 2592 2016 0 FreeSans 960 0 0 0 I18/VSS
flabel metal2 2592 4032 2592 4032 0 FreeSans 960 0 0 0 I18/VDD
flabel metal1 2562 3438 2622 3844 0 FreeSans 160 0 0 0 I18/MP0_IM0/D0
flabel metal1 2506 3276 2680 3348 0 FreeSans 160 0 0 0 I18/MP0_IM0/G0
flabel metal1 2706 3438 2766 3844 0 FreeSans 160 0 0 0 I18/MP0_IM0/S0
flabel metal1 2418 3438 2478 3844 0 FreeSans 160 0 0 0 I18/MP0_IM0/S1
flabel nwell 2732 3362 2756 3378 0 FreeSans 80 0 0 0 I18/MP0_IM0/BODY
flabel space 2304 3024 2448 4032 0 FreeSans 320 90 0 0 I18/MP0_IBNDR0/pmos_boundary
flabel space 2736 3024 2880 4032 0 FreeSans 320 90 0 0 I18/MP0_IBNDL0/pmos_boundary
flabel metal1 2706 2304 2766 2630 0 FreeSans 240 0 0 0 I18/MN0_IM0/S0
flabel metal1 2562 2304 2622 2630 0 FreeSans 240 0 0 0 I18/MN0_IM0/D0
flabel metal1 2418 2304 2478 2630 0 FreeSans 240 0 0 0 I18/MN0_IM0/S1
flabel metal1 2506 2700 2680 2772 0 FreeSans 240 0 0 0 I18/MN0_IM0/G0
rlabel pwell 2746 2670 2776 2692 1 I18/MN0_IM0/BODY
flabel space 2304 2016 2448 3024 0 FreeSans 320 90 0 0 I18/MN0_IBNDR0/nmos_boundary
flabel space 2736 2016 2880 3024 0 FreeSans 320 90 0 0 I18/MN0_IBNDL0/nmos_boundary
flabel metal3 3024 3024 3024 3024 0 FreeSans 480 90 0 0 I19/I
flabel metal3 3168 3024 3168 3024 0 FreeSans 480 90 0 0 I19/O
flabel metal2 3168 2016 3168 2016 0 FreeSans 960 0 0 0 I19/VSS
flabel metal2 3168 4032 3168 4032 0 FreeSans 960 0 0 0 I19/VDD
flabel metal1 3138 3438 3198 3844 0 FreeSans 160 0 0 0 I19/MP0_IM0/D0
flabel metal1 3080 3276 3254 3348 0 FreeSans 160 0 0 0 I19/MP0_IM0/G0
flabel metal1 2994 3438 3054 3844 0 FreeSans 160 0 0 0 I19/MP0_IM0/S0
flabel metal1 3282 3438 3342 3844 0 FreeSans 160 0 0 0 I19/MP0_IM0/S1
flabel nwell 3004 3362 3028 3378 0 FreeSans 80 0 0 0 I19/MP0_IM0/BODY
flabel space 3312 3024 3456 4032 0 FreeSans 320 90 0 0 I19/MP0_IBNDR0/pmos_boundary
flabel space 2880 3024 3024 4032 0 FreeSans 320 90 0 0 I19/MP0_IBNDL0/pmos_boundary
flabel metal1 2994 2304 3054 2630 0 FreeSans 240 0 0 0 I19/MN0_IM0/S0
flabel metal1 3138 2304 3198 2630 0 FreeSans 240 0 0 0 I19/MN0_IM0/D0
flabel metal1 3282 2304 3342 2630 0 FreeSans 240 0 0 0 I19/MN0_IM0/S1
flabel metal1 3080 2700 3254 2772 0 FreeSans 240 0 0 0 I19/MN0_IM0/G0
rlabel pwell 2984 2670 3014 2692 1 I19/MN0_IM0/BODY
flabel space 3312 2016 3456 3024 0 FreeSans 320 90 0 0 I19/MN0_IBNDR0/nmos_boundary
flabel space 2880 2016 3024 3024 0 FreeSans 320 90 0 0 I19/MN0_IBNDL0/nmos_boundary
flabel space 3888 3008 4032 4032 0 FreeSans 320 90 0 0 TAP1_1/MPT0_IBNDR0/ptap_boundary
flabel space 3456 3008 3600 4032 0 FreeSans 320 90 0 0 TAP1_1/MPT0_IBNDL0/ptap_boundary
flabel space 3888 2016 4032 3040 0 FreeSans 320 90 0 0 TAP1_1/MNT0_IBNDR0/ntap_boundary
flabel space 3456 2016 3600 3040 0 FreeSans 320 90 0 0 TAP1_1/MNT0_IBNDL0/ntap_boundary
flabel space 5616 0 5760 1024 0 FreeSans 320 90 0 0 TAP0_1/MPT0_IBNDR0/ptap_boundary
flabel space 5184 0 5328 1024 0 FreeSans 320 90 0 0 TAP0_1/MPT0_IBNDL0/ptap_boundary
flabel space 5616 992 5760 2016 0 FreeSans 320 90 0 0 TAP0_1/MNT0_IBNDR0/ntap_boundary
flabel space 5184 992 5328 2016 0 FreeSans 320 90 0 0 TAP0_1/MNT0_IBNDL0/ntap_boundary
flabel metal3 5472 3024 5472 3024 0 FreeSans 480 90 0 0 I20/I
flabel metal3 4176 3024 4176 3024 0 FreeSans 480 90 0 0 I20/CLK
flabel metal3 10368 3024 10368 3024 0 FreeSans 480 90 0 0 I20/O
flabel metal2 7344 2016 7344 2016 0 FreeSans 960 0 0 0 I20/VSS
flabel metal2 7344 4032 7344 4032 0 FreeSans 960 0 0 0 I20/VDD
flabel metal3 4176 3024 4176 3024 0 FreeSans 480 90 0 0 I20/inv0/I
flabel metal3 4320 3024 4320 3024 0 FreeSans 480 90 0 0 I20/inv0/O
flabel metal2 4320 2016 4320 2016 0 FreeSans 960 0 0 0 I20/inv0/VSS
flabel metal2 4320 4032 4320 4032 0 FreeSans 960 0 0 0 I20/inv0/VDD
flabel metal1 4290 3438 4350 3844 0 FreeSans 160 0 0 0 I20/inv0/MP0_IM0/D0
flabel metal1 4232 3276 4406 3348 0 FreeSans 160 0 0 0 I20/inv0/MP0_IM0/G0
flabel metal1 4146 3438 4206 3844 0 FreeSans 160 0 0 0 I20/inv0/MP0_IM0/S0
flabel metal1 4434 3438 4494 3844 0 FreeSans 160 0 0 0 I20/inv0/MP0_IM0/S1
flabel nwell 4156 3362 4180 3378 0 FreeSans 80 0 0 0 I20/inv0/MP0_IM0/BODY
flabel space 4464 3024 4608 4032 0 FreeSans 320 90 0 0 I20/inv0/MP0_IBNDR0/pmos_boundary
flabel space 4032 3024 4176 4032 0 FreeSans 320 90 0 0 I20/inv0/MP0_IBNDL0/pmos_boundary
flabel metal1 4146 2304 4206 2630 0 FreeSans 240 0 0 0 I20/inv0/MN0_IM0/S0
flabel metal1 4290 2304 4350 2630 0 FreeSans 240 0 0 0 I20/inv0/MN0_IM0/D0
flabel metal1 4434 2304 4494 2630 0 FreeSans 240 0 0 0 I20/inv0/MN0_IM0/S1
flabel metal1 4232 2700 4406 2772 0 FreeSans 240 0 0 0 I20/inv0/MN0_IM0/G0
rlabel pwell 4136 2670 4166 2692 1 I20/inv0/MN0_IM0/BODY
flabel space 4464 2016 4608 3024 0 FreeSans 320 90 0 0 I20/inv0/MN0_IBNDR0/nmos_boundary
flabel space 4032 2016 4176 3024 0 FreeSans 320 90 0 0 I20/inv0/MN0_IBNDL0/nmos_boundary
flabel metal3 4752 3024 4752 3024 0 FreeSans 480 90 0 0 I20/inv1/I
flabel metal3 4896 3024 4896 3024 0 FreeSans 480 90 0 0 I20/inv1/O
flabel metal2 4896 2016 4896 2016 0 FreeSans 960 0 0 0 I20/inv1/VSS
flabel metal2 4896 4032 4896 4032 0 FreeSans 960 0 0 0 I20/inv1/VDD
flabel metal1 4866 3438 4926 3844 0 FreeSans 160 0 0 0 I20/inv1/MP0_IM0/D0
flabel metal1 4808 3276 4982 3348 0 FreeSans 160 0 0 0 I20/inv1/MP0_IM0/G0
flabel metal1 4722 3438 4782 3844 0 FreeSans 160 0 0 0 I20/inv1/MP0_IM0/S0
flabel metal1 5010 3438 5070 3844 0 FreeSans 160 0 0 0 I20/inv1/MP0_IM0/S1
flabel nwell 4732 3362 4756 3378 0 FreeSans 80 0 0 0 I20/inv1/MP0_IM0/BODY
flabel space 5040 3024 5184 4032 0 FreeSans 320 90 0 0 I20/inv1/MP0_IBNDR0/pmos_boundary
flabel space 4608 3024 4752 4032 0 FreeSans 320 90 0 0 I20/inv1/MP0_IBNDL0/pmos_boundary
flabel metal1 4722 2304 4782 2630 0 FreeSans 240 0 0 0 I20/inv1/MN0_IM0/S0
flabel metal1 4866 2304 4926 2630 0 FreeSans 240 0 0 0 I20/inv1/MN0_IM0/D0
flabel metal1 5010 2304 5070 2630 0 FreeSans 240 0 0 0 I20/inv1/MN0_IM0/S1
flabel metal1 4808 2700 4982 2772 0 FreeSans 240 0 0 0 I20/inv1/MN0_IM0/G0
rlabel pwell 4712 2670 4742 2692 1 I20/inv1/MN0_IM0/BODY
flabel space 5040 2016 5184 3024 0 FreeSans 320 90 0 0 I20/inv1/MN0_IBNDR0/nmos_boundary
flabel space 4608 2016 4752 3024 0 FreeSans 320 90 0 0 I20/inv1/MN0_IBNDL0/nmos_boundary
flabel metal3 5472 3024 5472 3024 0 FreeSans 480 90 0 0 I20/tinv0/I
flabel metal3 6192 3024 6192 3024 0 FreeSans 480 90 0 0 I20/tinv0/EN
flabel metal3 5904 3024 5904 3024 0 FreeSans 480 90 0 0 I20/tinv0/ENB
flabel metal3 6048 3024 6048 3024 0 FreeSans 480 90 0 0 I20/tinv0/O
flabel metal2 5760 2016 5760 2016 0 FreeSans 960 0 0 0 I20/tinv0/VSS
flabel metal2 5760 4032 5760 4032 0 FreeSans 960 0 0 0 I20/tinv0/VDD
flabel metal1 6018 3438 6078 3844 0 FreeSans 160 0 0 0 I20/tinv0/MP1_IM0/D0
flabel metal1 5960 3276 6134 3348 0 FreeSans 160 0 0 0 I20/tinv0/MP1_IM0/G0
flabel metal1 5874 3438 5934 3844 0 FreeSans 160 0 0 0 I20/tinv0/MP1_IM0/S0
flabel metal1 6162 3438 6222 3844 0 FreeSans 160 0 0 0 I20/tinv0/MP1_IM0/S1
flabel nwell 5884 3362 5908 3378 0 FreeSans 80 0 0 0 I20/tinv0/MP1_IM0/BODY
flabel space 6192 3024 6336 4032 0 FreeSans 320 90 0 0 I20/tinv0/MP1_IBNDR0/pmos_boundary
flabel space 5760 3024 5904 4032 0 FreeSans 320 90 0 0 I20/tinv0/MP1_IBNDL0/pmos_boundary
flabel metal1 5442 3438 5502 3844 0 FreeSans 160 0 0 0 I20/tinv0/MP0_IM0/D0
flabel metal1 5384 3276 5558 3348 0 FreeSans 160 0 0 0 I20/tinv0/MP0_IM0/G0
flabel metal1 5298 3438 5358 3844 0 FreeSans 160 0 0 0 I20/tinv0/MP0_IM0/S0
flabel metal1 5586 3438 5646 3844 0 FreeSans 160 0 0 0 I20/tinv0/MP0_IM0/S1
flabel nwell 5308 3362 5332 3378 0 FreeSans 80 0 0 0 I20/tinv0/MP0_IM0/BODY
flabel space 5616 3024 5760 4032 0 FreeSans 320 90 0 0 I20/tinv0/MP0_IBNDR0/pmos_boundary
flabel space 5184 3024 5328 4032 0 FreeSans 320 90 0 0 I20/tinv0/MP0_IBNDL0/pmos_boundary
flabel metal1 5874 2304 5934 2630 0 FreeSans 240 0 0 0 I20/tinv0/MN1_IM0/S0
flabel metal1 6018 2304 6078 2630 0 FreeSans 240 0 0 0 I20/tinv0/MN1_IM0/D0
flabel metal1 6162 2304 6222 2630 0 FreeSans 240 0 0 0 I20/tinv0/MN1_IM0/S1
flabel metal1 5960 2700 6134 2772 0 FreeSans 240 0 0 0 I20/tinv0/MN1_IM0/G0
rlabel pwell 5864 2670 5894 2692 1 I20/tinv0/MN1_IM0/BODY
flabel space 6192 2016 6336 3024 0 FreeSans 320 90 0 0 I20/tinv0/MN1_IBNDR0/nmos_boundary
flabel space 5760 2016 5904 3024 0 FreeSans 320 90 0 0 I20/tinv0/MN1_IBNDL0/nmos_boundary
flabel metal1 5298 2304 5358 2630 0 FreeSans 240 0 0 0 I20/tinv0/MN0_IM0/S0
flabel metal1 5442 2304 5502 2630 0 FreeSans 240 0 0 0 I20/tinv0/MN0_IM0/D0
flabel metal1 5586 2304 5646 2630 0 FreeSans 240 0 0 0 I20/tinv0/MN0_IM0/S1
flabel metal1 5384 2700 5558 2772 0 FreeSans 240 0 0 0 I20/tinv0/MN0_IM0/G0
rlabel pwell 5288 2670 5318 2692 1 I20/tinv0/MN0_IM0/BODY
flabel space 5616 2016 5760 3024 0 FreeSans 320 90 0 0 I20/tinv0/MN0_IBNDR0/nmos_boundary
flabel space 5184 2016 5328 3024 0 FreeSans 320 90 0 0 I20/tinv0/MN0_IBNDL0/nmos_boundary
flabel metal3 6480 3024 6480 3024 0 FreeSans 480 90 0 0 I20/tinv_small0/I
flabel metal3 6768 3024 6768 3024 0 FreeSans 480 90 0 0 I20/tinv_small0/O
flabel metal3 6912 3024 6912 3024 0 FreeSans 480 90 0 0 I20/tinv_small0/EN
flabel metal3 6624 3024 6624 3024 0 FreeSans 480 90 0 0 I20/tinv_small0/ENB
flabel metal2 6768 2016 6768 2016 0 FreeSans 960 0 0 0 I20/tinv_small0/VSS
flabel metal2 6768 4032 6768 4032 0 FreeSans 960 0 0 0 I20/tinv_small0/VDD
flabel metal1 6446 3276 6536 3348 0 FreeSans 160 0 0 0 I20/tinv_small0/pstack/G0
flabel metal1 6710 3276 6800 3348 0 FreeSans 160 0 0 0 I20/tinv_small0/pstack/G1
flabel metal1 6450 3438 6510 3844 0 FreeSans 160 0 0 0 I20/tinv_small0/pstack/S0
flabel nwell 6460 3362 6484 3378 0 FreeSans 80 0 0 0 I20/tinv_small0/pstack/BODY
flabel metal1 6738 3438 6798 3844 0 FreeSans 160 0 0 0 I20/tinv_small0/pstack/D0
flabel space 7056 3024 7200 4032 0 FreeSans 320 90 0 0 I20/tinv_small0/pspace1/PMOS_SPACE
flabel space 6912 3024 7056 4032 0 FreeSans 320 90 0 0 I20/tinv_small0/pspace0/PMOS_SPACE
flabel space 6768 3024 6912 4032 0 FreeSans 320 90 0 0 I20/tinv_small0/pbndr/pmos_boundary
flabel space 6336 3024 6480 4032 0 FreeSans 320 90 0 0 I20/tinv_small0/pbndl/pmos_boundary
flabel metal1 6446 2700 6536 2772 0 FreeSans 160 0 0 0 I20/tinv_small0/nstack/G0
flabel metal1 6710 2700 6800 2772 0 FreeSans 160 0 0 0 I20/tinv_small0/nstack/G1
flabel metal1 6450 2304 6510 2630 0 FreeSans 160 0 0 0 I20/tinv_small0/nstack/S0
rlabel pwell 6440 2670 6470 2692 1 I20/tinv_small0/nstack/BODY
flabel metal1 6738 2304 6798 2630 0 FreeSans 160 0 0 0 I20/tinv_small0/nstack/D0
flabel space 7056 2016 7200 3024 0 FreeSans 320 90 0 0 I20/tinv_small0/nspace1/NMOS_SPACE
flabel space 6912 2016 7056 3024 0 FreeSans 320 90 0 0 I20/tinv_small0/nspace0/NMOS_SPACE
flabel space 6768 2016 6912 3024 0 FreeSans 320 90 0 0 I20/tinv_small0/nbndr/nmos_boundary
flabel space 6336 2016 6480 3024 0 FreeSans 320 90 0 0 I20/tinv_small0/nbndl/nmos_boundary
flabel space 6912 2016 7056 3040 0 FreeSans 320 90 0 0 I20/MNT0_IBNDL0/ntap_boundary
flabel space 6912 3008 7056 4032 0 FreeSans 320 90 0 0 I20/MPT0_IBNDL0/ptap_boundary
flabel space 7344 2016 7488 3040 0 FreeSans 320 90 0 0 I20/MNT0_IBNDR0/ntap_boundary
flabel space 7344 3008 7488 4032 0 FreeSans 320 90 0 0 I20/MPT0_IBNDR0/ptap_boundary
flabel metal3 7632 3024 7632 3024 0 FreeSans 480 90 0 0 I20/inv2/I
flabel metal3 7776 3024 7776 3024 0 FreeSans 480 90 0 0 I20/inv2/O
flabel metal2 7776 2016 7776 2016 0 FreeSans 960 0 0 0 I20/inv2/VSS
flabel metal2 7776 4032 7776 4032 0 FreeSans 960 0 0 0 I20/inv2/VDD
flabel metal1 7746 3438 7806 3844 0 FreeSans 160 0 0 0 I20/inv2/MP0_IM0/D0
flabel metal1 7688 3276 7862 3348 0 FreeSans 160 0 0 0 I20/inv2/MP0_IM0/G0
flabel metal1 7602 3438 7662 3844 0 FreeSans 160 0 0 0 I20/inv2/MP0_IM0/S0
flabel metal1 7890 3438 7950 3844 0 FreeSans 160 0 0 0 I20/inv2/MP0_IM0/S1
flabel nwell 7612 3362 7636 3378 0 FreeSans 80 0 0 0 I20/inv2/MP0_IM0/BODY
flabel space 7920 3024 8064 4032 0 FreeSans 320 90 0 0 I20/inv2/MP0_IBNDR0/pmos_boundary
flabel space 7488 3024 7632 4032 0 FreeSans 320 90 0 0 I20/inv2/MP0_IBNDL0/pmos_boundary
flabel metal1 7602 2304 7662 2630 0 FreeSans 240 0 0 0 I20/inv2/MN0_IM0/S0
flabel metal1 7746 2304 7806 2630 0 FreeSans 240 0 0 0 I20/inv2/MN0_IM0/D0
flabel metal1 7890 2304 7950 2630 0 FreeSans 240 0 0 0 I20/inv2/MN0_IM0/S1
flabel metal1 7688 2700 7862 2772 0 FreeSans 240 0 0 0 I20/inv2/MN0_IM0/G0
rlabel pwell 7592 2670 7622 2692 1 I20/inv2/MN0_IM0/BODY
flabel space 7920 2016 8064 3024 0 FreeSans 320 90 0 0 I20/inv2/MN0_IBNDR0/nmos_boundary
flabel space 7488 2016 7632 3024 0 FreeSans 320 90 0 0 I20/inv2/MN0_IBNDL0/nmos_boundary
flabel metal3 8352 3024 8352 3024 0 FreeSans 480 90 0 0 I20/tinv1/I
flabel metal3 9072 3024 9072 3024 0 FreeSans 480 90 0 0 I20/tinv1/EN
flabel metal3 8784 3024 8784 3024 0 FreeSans 480 90 0 0 I20/tinv1/ENB
flabel metal3 8928 3024 8928 3024 0 FreeSans 480 90 0 0 I20/tinv1/O
flabel metal2 8640 2016 8640 2016 0 FreeSans 960 0 0 0 I20/tinv1/VSS
flabel metal2 8640 4032 8640 4032 0 FreeSans 960 0 0 0 I20/tinv1/VDD
flabel metal1 8898 3438 8958 3844 0 FreeSans 160 0 0 0 I20/tinv1/MP1_IM0/D0
flabel metal1 8840 3276 9014 3348 0 FreeSans 160 0 0 0 I20/tinv1/MP1_IM0/G0
flabel metal1 8754 3438 8814 3844 0 FreeSans 160 0 0 0 I20/tinv1/MP1_IM0/S0
flabel metal1 9042 3438 9102 3844 0 FreeSans 160 0 0 0 I20/tinv1/MP1_IM0/S1
flabel nwell 8764 3362 8788 3378 0 FreeSans 80 0 0 0 I20/tinv1/MP1_IM0/BODY
flabel space 9072 3024 9216 4032 0 FreeSans 320 90 0 0 I20/tinv1/MP1_IBNDR0/pmos_boundary
flabel space 8640 3024 8784 4032 0 FreeSans 320 90 0 0 I20/tinv1/MP1_IBNDL0/pmos_boundary
flabel metal1 8322 3438 8382 3844 0 FreeSans 160 0 0 0 I20/tinv1/MP0_IM0/D0
flabel metal1 8264 3276 8438 3348 0 FreeSans 160 0 0 0 I20/tinv1/MP0_IM0/G0
flabel metal1 8178 3438 8238 3844 0 FreeSans 160 0 0 0 I20/tinv1/MP0_IM0/S0
flabel metal1 8466 3438 8526 3844 0 FreeSans 160 0 0 0 I20/tinv1/MP0_IM0/S1
flabel nwell 8188 3362 8212 3378 0 FreeSans 80 0 0 0 I20/tinv1/MP0_IM0/BODY
flabel space 8496 3024 8640 4032 0 FreeSans 320 90 0 0 I20/tinv1/MP0_IBNDR0/pmos_boundary
flabel space 8064 3024 8208 4032 0 FreeSans 320 90 0 0 I20/tinv1/MP0_IBNDL0/pmos_boundary
flabel metal1 8754 2304 8814 2630 0 FreeSans 240 0 0 0 I20/tinv1/MN1_IM0/S0
flabel metal1 8898 2304 8958 2630 0 FreeSans 240 0 0 0 I20/tinv1/MN1_IM0/D0
flabel metal1 9042 2304 9102 2630 0 FreeSans 240 0 0 0 I20/tinv1/MN1_IM0/S1
flabel metal1 8840 2700 9014 2772 0 FreeSans 240 0 0 0 I20/tinv1/MN1_IM0/G0
rlabel pwell 8744 2670 8774 2692 1 I20/tinv1/MN1_IM0/BODY
flabel space 9072 2016 9216 3024 0 FreeSans 320 90 0 0 I20/tinv1/MN1_IBNDR0/nmos_boundary
flabel space 8640 2016 8784 3024 0 FreeSans 320 90 0 0 I20/tinv1/MN1_IBNDL0/nmos_boundary
flabel metal1 8178 2304 8238 2630 0 FreeSans 240 0 0 0 I20/tinv1/MN0_IM0/S0
flabel metal1 8322 2304 8382 2630 0 FreeSans 240 0 0 0 I20/tinv1/MN0_IM0/D0
flabel metal1 8466 2304 8526 2630 0 FreeSans 240 0 0 0 I20/tinv1/MN0_IM0/S1
flabel metal1 8264 2700 8438 2772 0 FreeSans 240 0 0 0 I20/tinv1/MN0_IM0/G0
rlabel pwell 8168 2670 8198 2692 1 I20/tinv1/MN0_IM0/BODY
flabel space 8496 2016 8640 3024 0 FreeSans 320 90 0 0 I20/tinv1/MN0_IBNDR0/nmos_boundary
flabel space 8064 2016 8208 3024 0 FreeSans 320 90 0 0 I20/tinv1/MN0_IBNDL0/nmos_boundary
flabel metal3 10224 3024 10224 3024 0 FreeSans 480 90 0 0 I20/inv3/I
flabel metal3 10368 3024 10368 3024 0 FreeSans 480 90 0 0 I20/inv3/O
flabel metal2 10368 2016 10368 2016 0 FreeSans 960 0 0 0 I20/inv3/VSS
flabel metal2 10368 4032 10368 4032 0 FreeSans 960 0 0 0 I20/inv3/VDD
flabel metal1 10338 3438 10398 3844 0 FreeSans 160 0 0 0 I20/inv3/MP0_IM0/D0
flabel metal1 10280 3276 10454 3348 0 FreeSans 160 0 0 0 I20/inv3/MP0_IM0/G0
flabel metal1 10194 3438 10254 3844 0 FreeSans 160 0 0 0 I20/inv3/MP0_IM0/S0
flabel metal1 10482 3438 10542 3844 0 FreeSans 160 0 0 0 I20/inv3/MP0_IM0/S1
flabel nwell 10204 3362 10228 3378 0 FreeSans 80 0 0 0 I20/inv3/MP0_IM0/BODY
flabel space 10512 3024 10656 4032 0 FreeSans 320 90 0 0 I20/inv3/MP0_IBNDR0/pmos_boundary
flabel space 10080 3024 10224 4032 0 FreeSans 320 90 0 0 I20/inv3/MP0_IBNDL0/pmos_boundary
flabel metal1 10194 2304 10254 2630 0 FreeSans 240 0 0 0 I20/inv3/MN0_IM0/S0
flabel metal1 10338 2304 10398 2630 0 FreeSans 240 0 0 0 I20/inv3/MN0_IM0/D0
flabel metal1 10482 2304 10542 2630 0 FreeSans 240 0 0 0 I20/inv3/MN0_IM0/S1
flabel metal1 10280 2700 10454 2772 0 FreeSans 240 0 0 0 I20/inv3/MN0_IM0/G0
rlabel pwell 10184 2670 10214 2692 1 I20/inv3/MN0_IM0/BODY
flabel space 10512 2016 10656 3024 0 FreeSans 320 90 0 0 I20/inv3/MN0_IBNDR0/nmos_boundary
flabel space 10080 2016 10224 3024 0 FreeSans 320 90 0 0 I20/inv3/MN0_IBNDL0/nmos_boundary
flabel metal3 9360 3024 9360 3024 0 FreeSans 480 90 0 0 I20/tinv_small1/I
flabel metal3 9648 3024 9648 3024 0 FreeSans 480 90 0 0 I20/tinv_small1/O
flabel metal3 9792 3024 9792 3024 0 FreeSans 480 90 0 0 I20/tinv_small1/EN
flabel metal3 9504 3024 9504 3024 0 FreeSans 480 90 0 0 I20/tinv_small1/ENB
flabel metal2 9648 2016 9648 2016 0 FreeSans 960 0 0 0 I20/tinv_small1/VSS
flabel metal2 9648 4032 9648 4032 0 FreeSans 960 0 0 0 I20/tinv_small1/VDD
flabel metal1 9326 3276 9416 3348 0 FreeSans 160 0 0 0 I20/tinv_small1/pstack/G0
flabel metal1 9590 3276 9680 3348 0 FreeSans 160 0 0 0 I20/tinv_small1/pstack/G1
flabel metal1 9330 3438 9390 3844 0 FreeSans 160 0 0 0 I20/tinv_small1/pstack/S0
flabel nwell 9340 3362 9364 3378 0 FreeSans 80 0 0 0 I20/tinv_small1/pstack/BODY
flabel metal1 9618 3438 9678 3844 0 FreeSans 160 0 0 0 I20/tinv_small1/pstack/D0
flabel space 9936 3024 10080 4032 0 FreeSans 320 90 0 0 I20/tinv_small1/pspace1/PMOS_SPACE
flabel space 9792 3024 9936 4032 0 FreeSans 320 90 0 0 I20/tinv_small1/pspace0/PMOS_SPACE
flabel space 9648 3024 9792 4032 0 FreeSans 320 90 0 0 I20/tinv_small1/pbndr/pmos_boundary
flabel space 9216 3024 9360 4032 0 FreeSans 320 90 0 0 I20/tinv_small1/pbndl/pmos_boundary
flabel metal1 9326 2700 9416 2772 0 FreeSans 160 0 0 0 I20/tinv_small1/nstack/G0
flabel metal1 9590 2700 9680 2772 0 FreeSans 160 0 0 0 I20/tinv_small1/nstack/G1
flabel metal1 9330 2304 9390 2630 0 FreeSans 160 0 0 0 I20/tinv_small1/nstack/S0
rlabel pwell 9320 2670 9350 2692 1 I20/tinv_small1/nstack/BODY
flabel metal1 9618 2304 9678 2630 0 FreeSans 160 0 0 0 I20/tinv_small1/nstack/D0
flabel space 9936 2016 10080 3024 0 FreeSans 320 90 0 0 I20/tinv_small1/nspace1/NMOS_SPACE
flabel space 9792 2016 9936 3024 0 FreeSans 320 90 0 0 I20/tinv_small1/nspace0/NMOS_SPACE
flabel space 9648 2016 9792 3024 0 FreeSans 320 90 0 0 I20/tinv_small1/nbndr/nmos_boundary
flabel space 9216 2016 9360 3024 0 FreeSans 320 90 0 0 I20/tinv_small1/nbndl/nmos_boundary
flabel metal3 7200 1008 7200 1008 0 FreeSans 480 90 0 0 I2/I
flabel metal3 5904 1008 5904 1008 0 FreeSans 480 90 0 0 I2/CLK
flabel metal3 12096 1008 12096 1008 0 FreeSans 480 90 0 0 I2/O
flabel metal2 9072 2016 9072 2016 0 FreeSans 960 0 0 0 I2/VSS
flabel metal2 9072 0 9072 0 0 FreeSans 960 0 0 0 I2/VDD
flabel metal3 5904 1008 5904 1008 0 FreeSans 480 90 0 0 I2/inv0/I
flabel metal3 6048 1008 6048 1008 0 FreeSans 480 90 0 0 I2/inv0/O
flabel metal2 6048 2016 6048 2016 0 FreeSans 960 0 0 0 I2/inv0/VSS
flabel metal2 6048 0 6048 0 0 FreeSans 960 0 0 0 I2/inv0/VDD
flabel metal1 6018 188 6078 594 0 FreeSans 160 0 0 0 I2/inv0/MP0_IM0/D0
flabel metal1 5960 684 6134 756 0 FreeSans 160 0 0 0 I2/inv0/MP0_IM0/G0
flabel metal1 5874 188 5934 594 0 FreeSans 160 0 0 0 I2/inv0/MP0_IM0/S0
flabel metal1 6162 188 6222 594 0 FreeSans 160 0 0 0 I2/inv0/MP0_IM0/S1
flabel nwell 5884 654 5908 670 0 FreeSans 80 0 0 0 I2/inv0/MP0_IM0/BODY
flabel space 6192 0 6336 1008 0 FreeSans 320 90 0 0 I2/inv0/MP0_IBNDR0/pmos_boundary
flabel space 5760 0 5904 1008 0 FreeSans 320 90 0 0 I2/inv0/MP0_IBNDL0/pmos_boundary
flabel metal1 5874 1402 5934 1728 0 FreeSans 240 0 0 0 I2/inv0/MN0_IM0/S0
flabel metal1 6018 1402 6078 1728 0 FreeSans 240 0 0 0 I2/inv0/MN0_IM0/D0
flabel metal1 6162 1402 6222 1728 0 FreeSans 240 0 0 0 I2/inv0/MN0_IM0/S1
flabel metal1 5960 1260 6134 1332 0 FreeSans 240 0 0 0 I2/inv0/MN0_IM0/G0
rlabel pwell 5864 1340 5894 1362 5 I2/inv0/MN0_IM0/BODY
flabel space 6192 1008 6336 2016 0 FreeSans 320 90 0 0 I2/inv0/MN0_IBNDR0/nmos_boundary
flabel space 5760 1008 5904 2016 0 FreeSans 320 90 0 0 I2/inv0/MN0_IBNDL0/nmos_boundary
flabel metal3 6480 1008 6480 1008 0 FreeSans 480 90 0 0 I2/inv1/I
flabel metal3 6624 1008 6624 1008 0 FreeSans 480 90 0 0 I2/inv1/O
flabel metal2 6624 2016 6624 2016 0 FreeSans 960 0 0 0 I2/inv1/VSS
flabel metal2 6624 0 6624 0 0 FreeSans 960 0 0 0 I2/inv1/VDD
flabel metal1 6594 188 6654 594 0 FreeSans 160 0 0 0 I2/inv1/MP0_IM0/D0
flabel metal1 6536 684 6710 756 0 FreeSans 160 0 0 0 I2/inv1/MP0_IM0/G0
flabel metal1 6450 188 6510 594 0 FreeSans 160 0 0 0 I2/inv1/MP0_IM0/S0
flabel metal1 6738 188 6798 594 0 FreeSans 160 0 0 0 I2/inv1/MP0_IM0/S1
flabel nwell 6460 654 6484 670 0 FreeSans 80 0 0 0 I2/inv1/MP0_IM0/BODY
flabel space 6768 0 6912 1008 0 FreeSans 320 90 0 0 I2/inv1/MP0_IBNDR0/pmos_boundary
flabel space 6336 0 6480 1008 0 FreeSans 320 90 0 0 I2/inv1/MP0_IBNDL0/pmos_boundary
flabel metal1 6450 1402 6510 1728 0 FreeSans 240 0 0 0 I2/inv1/MN0_IM0/S0
flabel metal1 6594 1402 6654 1728 0 FreeSans 240 0 0 0 I2/inv1/MN0_IM0/D0
flabel metal1 6738 1402 6798 1728 0 FreeSans 240 0 0 0 I2/inv1/MN0_IM0/S1
flabel metal1 6536 1260 6710 1332 0 FreeSans 240 0 0 0 I2/inv1/MN0_IM0/G0
rlabel pwell 6440 1340 6470 1362 5 I2/inv1/MN0_IM0/BODY
flabel space 6768 1008 6912 2016 0 FreeSans 320 90 0 0 I2/inv1/MN0_IBNDR0/nmos_boundary
flabel space 6336 1008 6480 2016 0 FreeSans 320 90 0 0 I2/inv1/MN0_IBNDL0/nmos_boundary
flabel metal3 7200 1008 7200 1008 0 FreeSans 480 90 0 0 I2/tinv0/I
flabel metal3 7920 1008 7920 1008 0 FreeSans 480 90 0 0 I2/tinv0/EN
flabel metal3 7632 1008 7632 1008 0 FreeSans 480 90 0 0 I2/tinv0/ENB
flabel metal3 7776 1008 7776 1008 0 FreeSans 480 90 0 0 I2/tinv0/O
flabel metal2 7488 2016 7488 2016 0 FreeSans 960 0 0 0 I2/tinv0/VSS
flabel metal2 7488 0 7488 0 0 FreeSans 960 0 0 0 I2/tinv0/VDD
flabel metal1 7746 188 7806 594 0 FreeSans 160 0 0 0 I2/tinv0/MP1_IM0/D0
flabel metal1 7688 684 7862 756 0 FreeSans 160 0 0 0 I2/tinv0/MP1_IM0/G0
flabel metal1 7602 188 7662 594 0 FreeSans 160 0 0 0 I2/tinv0/MP1_IM0/S0
flabel metal1 7890 188 7950 594 0 FreeSans 160 0 0 0 I2/tinv0/MP1_IM0/S1
flabel nwell 7612 654 7636 670 0 FreeSans 80 0 0 0 I2/tinv0/MP1_IM0/BODY
flabel space 7920 0 8064 1008 0 FreeSans 320 90 0 0 I2/tinv0/MP1_IBNDR0/pmos_boundary
flabel space 7488 0 7632 1008 0 FreeSans 320 90 0 0 I2/tinv0/MP1_IBNDL0/pmos_boundary
flabel metal1 7170 188 7230 594 0 FreeSans 160 0 0 0 I2/tinv0/MP0_IM0/D0
flabel metal1 7112 684 7286 756 0 FreeSans 160 0 0 0 I2/tinv0/MP0_IM0/G0
flabel metal1 7026 188 7086 594 0 FreeSans 160 0 0 0 I2/tinv0/MP0_IM0/S0
flabel metal1 7314 188 7374 594 0 FreeSans 160 0 0 0 I2/tinv0/MP0_IM0/S1
flabel nwell 7036 654 7060 670 0 FreeSans 80 0 0 0 I2/tinv0/MP0_IM0/BODY
flabel space 7344 0 7488 1008 0 FreeSans 320 90 0 0 I2/tinv0/MP0_IBNDR0/pmos_boundary
flabel space 6912 0 7056 1008 0 FreeSans 320 90 0 0 I2/tinv0/MP0_IBNDL0/pmos_boundary
flabel metal1 7602 1402 7662 1728 0 FreeSans 240 0 0 0 I2/tinv0/MN1_IM0/S0
flabel metal1 7746 1402 7806 1728 0 FreeSans 240 0 0 0 I2/tinv0/MN1_IM0/D0
flabel metal1 7890 1402 7950 1728 0 FreeSans 240 0 0 0 I2/tinv0/MN1_IM0/S1
flabel metal1 7688 1260 7862 1332 0 FreeSans 240 0 0 0 I2/tinv0/MN1_IM0/G0
rlabel pwell 7592 1340 7622 1362 5 I2/tinv0/MN1_IM0/BODY
flabel space 7920 1008 8064 2016 0 FreeSans 320 90 0 0 I2/tinv0/MN1_IBNDR0/nmos_boundary
flabel space 7488 1008 7632 2016 0 FreeSans 320 90 0 0 I2/tinv0/MN1_IBNDL0/nmos_boundary
flabel metal1 7026 1402 7086 1728 0 FreeSans 240 0 0 0 I2/tinv0/MN0_IM0/S0
flabel metal1 7170 1402 7230 1728 0 FreeSans 240 0 0 0 I2/tinv0/MN0_IM0/D0
flabel metal1 7314 1402 7374 1728 0 FreeSans 240 0 0 0 I2/tinv0/MN0_IM0/S1
flabel metal1 7112 1260 7286 1332 0 FreeSans 240 0 0 0 I2/tinv0/MN0_IM0/G0
rlabel pwell 7016 1340 7046 1362 5 I2/tinv0/MN0_IM0/BODY
flabel space 7344 1008 7488 2016 0 FreeSans 320 90 0 0 I2/tinv0/MN0_IBNDR0/nmos_boundary
flabel space 6912 1008 7056 2016 0 FreeSans 320 90 0 0 I2/tinv0/MN0_IBNDL0/nmos_boundary
flabel metal3 8208 1008 8208 1008 0 FreeSans 480 90 0 0 I2/tinv_small0/I
flabel metal3 8496 1008 8496 1008 0 FreeSans 480 90 0 0 I2/tinv_small0/O
flabel metal3 8640 1008 8640 1008 0 FreeSans 480 90 0 0 I2/tinv_small0/EN
flabel metal3 8352 1008 8352 1008 0 FreeSans 480 90 0 0 I2/tinv_small0/ENB
flabel metal2 8496 2016 8496 2016 0 FreeSans 960 0 0 0 I2/tinv_small0/VSS
flabel metal2 8496 0 8496 0 0 FreeSans 960 0 0 0 I2/tinv_small0/VDD
flabel metal1 8174 684 8264 756 0 FreeSans 160 0 0 0 I2/tinv_small0/pstack/G0
flabel metal1 8438 684 8528 756 0 FreeSans 160 0 0 0 I2/tinv_small0/pstack/G1
flabel metal1 8178 188 8238 594 0 FreeSans 160 0 0 0 I2/tinv_small0/pstack/S0
flabel nwell 8188 654 8212 670 0 FreeSans 80 0 0 0 I2/tinv_small0/pstack/BODY
flabel metal1 8466 188 8526 594 0 FreeSans 160 0 0 0 I2/tinv_small0/pstack/D0
flabel space 8784 0 8928 1008 0 FreeSans 320 90 0 0 I2/tinv_small0/pspace1/PMOS_SPACE
flabel space 8640 0 8784 1008 0 FreeSans 320 90 0 0 I2/tinv_small0/pspace0/PMOS_SPACE
flabel space 8496 0 8640 1008 0 FreeSans 320 90 0 0 I2/tinv_small0/pbndr/pmos_boundary
flabel space 8064 0 8208 1008 0 FreeSans 320 90 0 0 I2/tinv_small0/pbndl/pmos_boundary
flabel metal1 8174 1260 8264 1332 0 FreeSans 160 0 0 0 I2/tinv_small0/nstack/G0
flabel metal1 8438 1260 8528 1332 0 FreeSans 160 0 0 0 I2/tinv_small0/nstack/G1
flabel metal1 8178 1402 8238 1728 0 FreeSans 160 0 0 0 I2/tinv_small0/nstack/S0
rlabel pwell 8168 1340 8198 1362 5 I2/tinv_small0/nstack/BODY
flabel metal1 8466 1402 8526 1728 0 FreeSans 160 0 0 0 I2/tinv_small0/nstack/D0
flabel space 8784 1008 8928 2016 0 FreeSans 320 90 0 0 I2/tinv_small0/nspace1/NMOS_SPACE
flabel space 8640 1008 8784 2016 0 FreeSans 320 90 0 0 I2/tinv_small0/nspace0/NMOS_SPACE
flabel space 8496 1008 8640 2016 0 FreeSans 320 90 0 0 I2/tinv_small0/nbndr/nmos_boundary
flabel space 8064 1008 8208 2016 0 FreeSans 320 90 0 0 I2/tinv_small0/nbndl/nmos_boundary
flabel space 8640 992 8784 2016 0 FreeSans 320 90 0 0 I2/MNT0_IBNDL0/ntap_boundary
flabel space 8640 0 8784 1024 0 FreeSans 320 90 0 0 I2/MPT0_IBNDL0/ptap_boundary
flabel space 9072 992 9216 2016 0 FreeSans 320 90 0 0 I2/MNT0_IBNDR0/ntap_boundary
flabel space 9072 0 9216 1024 0 FreeSans 320 90 0 0 I2/MPT0_IBNDR0/ptap_boundary
flabel metal3 9360 1008 9360 1008 0 FreeSans 480 90 0 0 I2/inv2/I
flabel metal3 9504 1008 9504 1008 0 FreeSans 480 90 0 0 I2/inv2/O
flabel metal2 9504 2016 9504 2016 0 FreeSans 960 0 0 0 I2/inv2/VSS
flabel metal2 9504 0 9504 0 0 FreeSans 960 0 0 0 I2/inv2/VDD
flabel metal1 9474 188 9534 594 0 FreeSans 160 0 0 0 I2/inv2/MP0_IM0/D0
flabel metal1 9416 684 9590 756 0 FreeSans 160 0 0 0 I2/inv2/MP0_IM0/G0
flabel metal1 9330 188 9390 594 0 FreeSans 160 0 0 0 I2/inv2/MP0_IM0/S0
flabel metal1 9618 188 9678 594 0 FreeSans 160 0 0 0 I2/inv2/MP0_IM0/S1
flabel nwell 9340 654 9364 670 0 FreeSans 80 0 0 0 I2/inv2/MP0_IM0/BODY
flabel space 9648 0 9792 1008 0 FreeSans 320 90 0 0 I2/inv2/MP0_IBNDR0/pmos_boundary
flabel space 9216 0 9360 1008 0 FreeSans 320 90 0 0 I2/inv2/MP0_IBNDL0/pmos_boundary
flabel metal1 9330 1402 9390 1728 0 FreeSans 240 0 0 0 I2/inv2/MN0_IM0/S0
flabel metal1 9474 1402 9534 1728 0 FreeSans 240 0 0 0 I2/inv2/MN0_IM0/D0
flabel metal1 9618 1402 9678 1728 0 FreeSans 240 0 0 0 I2/inv2/MN0_IM0/S1
flabel metal1 9416 1260 9590 1332 0 FreeSans 240 0 0 0 I2/inv2/MN0_IM0/G0
rlabel pwell 9320 1340 9350 1362 5 I2/inv2/MN0_IM0/BODY
flabel space 9648 1008 9792 2016 0 FreeSans 320 90 0 0 I2/inv2/MN0_IBNDR0/nmos_boundary
flabel space 9216 1008 9360 2016 0 FreeSans 320 90 0 0 I2/inv2/MN0_IBNDL0/nmos_boundary
flabel metal3 10080 1008 10080 1008 0 FreeSans 480 90 0 0 I2/tinv1/I
flabel metal3 10800 1008 10800 1008 0 FreeSans 480 90 0 0 I2/tinv1/EN
flabel metal3 10512 1008 10512 1008 0 FreeSans 480 90 0 0 I2/tinv1/ENB
flabel metal3 10656 1008 10656 1008 0 FreeSans 480 90 0 0 I2/tinv1/O
flabel metal2 10368 2016 10368 2016 0 FreeSans 960 0 0 0 I2/tinv1/VSS
flabel metal2 10368 0 10368 0 0 FreeSans 960 0 0 0 I2/tinv1/VDD
flabel metal1 10626 188 10686 594 0 FreeSans 160 0 0 0 I2/tinv1/MP1_IM0/D0
flabel metal1 10568 684 10742 756 0 FreeSans 160 0 0 0 I2/tinv1/MP1_IM0/G0
flabel metal1 10482 188 10542 594 0 FreeSans 160 0 0 0 I2/tinv1/MP1_IM0/S0
flabel metal1 10770 188 10830 594 0 FreeSans 160 0 0 0 I2/tinv1/MP1_IM0/S1
flabel nwell 10492 654 10516 670 0 FreeSans 80 0 0 0 I2/tinv1/MP1_IM0/BODY
flabel space 10800 0 10944 1008 0 FreeSans 320 90 0 0 I2/tinv1/MP1_IBNDR0/pmos_boundary
flabel space 10368 0 10512 1008 0 FreeSans 320 90 0 0 I2/tinv1/MP1_IBNDL0/pmos_boundary
flabel metal1 10050 188 10110 594 0 FreeSans 160 0 0 0 I2/tinv1/MP0_IM0/D0
flabel metal1 9992 684 10166 756 0 FreeSans 160 0 0 0 I2/tinv1/MP0_IM0/G0
flabel metal1 9906 188 9966 594 0 FreeSans 160 0 0 0 I2/tinv1/MP0_IM0/S0
flabel metal1 10194 188 10254 594 0 FreeSans 160 0 0 0 I2/tinv1/MP0_IM0/S1
flabel nwell 9916 654 9940 670 0 FreeSans 80 0 0 0 I2/tinv1/MP0_IM0/BODY
flabel space 10224 0 10368 1008 0 FreeSans 320 90 0 0 I2/tinv1/MP0_IBNDR0/pmos_boundary
flabel space 9792 0 9936 1008 0 FreeSans 320 90 0 0 I2/tinv1/MP0_IBNDL0/pmos_boundary
flabel metal1 10482 1402 10542 1728 0 FreeSans 240 0 0 0 I2/tinv1/MN1_IM0/S0
flabel metal1 10626 1402 10686 1728 0 FreeSans 240 0 0 0 I2/tinv1/MN1_IM0/D0
flabel metal1 10770 1402 10830 1728 0 FreeSans 240 0 0 0 I2/tinv1/MN1_IM0/S1
flabel metal1 10568 1260 10742 1332 0 FreeSans 240 0 0 0 I2/tinv1/MN1_IM0/G0
rlabel pwell 10472 1340 10502 1362 5 I2/tinv1/MN1_IM0/BODY
flabel space 10800 1008 10944 2016 0 FreeSans 320 90 0 0 I2/tinv1/MN1_IBNDR0/nmos_boundary
flabel space 10368 1008 10512 2016 0 FreeSans 320 90 0 0 I2/tinv1/MN1_IBNDL0/nmos_boundary
flabel metal1 9906 1402 9966 1728 0 FreeSans 240 0 0 0 I2/tinv1/MN0_IM0/S0
flabel metal1 10050 1402 10110 1728 0 FreeSans 240 0 0 0 I2/tinv1/MN0_IM0/D0
flabel metal1 10194 1402 10254 1728 0 FreeSans 240 0 0 0 I2/tinv1/MN0_IM0/S1
flabel metal1 9992 1260 10166 1332 0 FreeSans 240 0 0 0 I2/tinv1/MN0_IM0/G0
rlabel pwell 9896 1340 9926 1362 5 I2/tinv1/MN0_IM0/BODY
flabel space 10224 1008 10368 2016 0 FreeSans 320 90 0 0 I2/tinv1/MN0_IBNDR0/nmos_boundary
flabel space 9792 1008 9936 2016 0 FreeSans 320 90 0 0 I2/tinv1/MN0_IBNDL0/nmos_boundary
flabel metal3 11952 1008 11952 1008 0 FreeSans 480 90 0 0 I2/inv3/I
flabel metal3 12096 1008 12096 1008 0 FreeSans 480 90 0 0 I2/inv3/O
flabel metal2 12096 2016 12096 2016 0 FreeSans 960 0 0 0 I2/inv3/VSS
flabel metal2 12096 0 12096 0 0 FreeSans 960 0 0 0 I2/inv3/VDD
flabel metal1 12066 188 12126 594 0 FreeSans 160 0 0 0 I2/inv3/MP0_IM0/D0
flabel metal1 12008 684 12182 756 0 FreeSans 160 0 0 0 I2/inv3/MP0_IM0/G0
flabel metal1 11922 188 11982 594 0 FreeSans 160 0 0 0 I2/inv3/MP0_IM0/S0
flabel metal1 12210 188 12270 594 0 FreeSans 160 0 0 0 I2/inv3/MP0_IM0/S1
flabel nwell 11932 654 11956 670 0 FreeSans 80 0 0 0 I2/inv3/MP0_IM0/BODY
flabel space 12240 0 12384 1008 0 FreeSans 320 90 0 0 I2/inv3/MP0_IBNDR0/pmos_boundary
flabel space 11808 0 11952 1008 0 FreeSans 320 90 0 0 I2/inv3/MP0_IBNDL0/pmos_boundary
flabel metal1 11922 1402 11982 1728 0 FreeSans 240 0 0 0 I2/inv3/MN0_IM0/S0
flabel metal1 12066 1402 12126 1728 0 FreeSans 240 0 0 0 I2/inv3/MN0_IM0/D0
flabel metal1 12210 1402 12270 1728 0 FreeSans 240 0 0 0 I2/inv3/MN0_IM0/S1
flabel metal1 12008 1260 12182 1332 0 FreeSans 240 0 0 0 I2/inv3/MN0_IM0/G0
rlabel pwell 11912 1340 11942 1362 5 I2/inv3/MN0_IM0/BODY
flabel space 12240 1008 12384 2016 0 FreeSans 320 90 0 0 I2/inv3/MN0_IBNDR0/nmos_boundary
flabel space 11808 1008 11952 2016 0 FreeSans 320 90 0 0 I2/inv3/MN0_IBNDL0/nmos_boundary
flabel metal3 11088 1008 11088 1008 0 FreeSans 480 90 0 0 I2/tinv_small1/I
flabel metal3 11376 1008 11376 1008 0 FreeSans 480 90 0 0 I2/tinv_small1/O
flabel metal3 11520 1008 11520 1008 0 FreeSans 480 90 0 0 I2/tinv_small1/EN
flabel metal3 11232 1008 11232 1008 0 FreeSans 480 90 0 0 I2/tinv_small1/ENB
flabel metal2 11376 2016 11376 2016 0 FreeSans 960 0 0 0 I2/tinv_small1/VSS
flabel metal2 11376 0 11376 0 0 FreeSans 960 0 0 0 I2/tinv_small1/VDD
flabel metal1 11054 684 11144 756 0 FreeSans 160 0 0 0 I2/tinv_small1/pstack/G0
flabel metal1 11318 684 11408 756 0 FreeSans 160 0 0 0 I2/tinv_small1/pstack/G1
flabel metal1 11058 188 11118 594 0 FreeSans 160 0 0 0 I2/tinv_small1/pstack/S0
flabel nwell 11068 654 11092 670 0 FreeSans 80 0 0 0 I2/tinv_small1/pstack/BODY
flabel metal1 11346 188 11406 594 0 FreeSans 160 0 0 0 I2/tinv_small1/pstack/D0
flabel space 11664 0 11808 1008 0 FreeSans 320 90 0 0 I2/tinv_small1/pspace1/PMOS_SPACE
flabel space 11520 0 11664 1008 0 FreeSans 320 90 0 0 I2/tinv_small1/pspace0/PMOS_SPACE
flabel space 11376 0 11520 1008 0 FreeSans 320 90 0 0 I2/tinv_small1/pbndr/pmos_boundary
flabel space 10944 0 11088 1008 0 FreeSans 320 90 0 0 I2/tinv_small1/pbndl/pmos_boundary
flabel metal1 11054 1260 11144 1332 0 FreeSans 160 0 0 0 I2/tinv_small1/nstack/G0
flabel metal1 11318 1260 11408 1332 0 FreeSans 160 0 0 0 I2/tinv_small1/nstack/G1
flabel metal1 11058 1402 11118 1728 0 FreeSans 160 0 0 0 I2/tinv_small1/nstack/S0
rlabel pwell 11048 1340 11078 1362 5 I2/tinv_small1/nstack/BODY
flabel metal1 11346 1402 11406 1728 0 FreeSans 160 0 0 0 I2/tinv_small1/nstack/D0
flabel space 11664 1008 11808 2016 0 FreeSans 320 90 0 0 I2/tinv_small1/nspace1/NMOS_SPACE
flabel space 11520 1008 11664 2016 0 FreeSans 320 90 0 0 I2/tinv_small1/nspace0/NMOS_SPACE
flabel space 11376 1008 11520 2016 0 FreeSans 320 90 0 0 I2/tinv_small1/nbndr/nmos_boundary
flabel space 10944 1008 11088 2016 0 FreeSans 320 90 0 0 I2/tinv_small1/nbndl/nmos_boundary
flabel metal3 1440 1008 1440 1008 0 FreeSans 480 90 0 0 I1/I0
flabel metal3 3744 1008 3744 1008 0 FreeSans 480 90 0 0 I1/I1
flabel metal3 2592 1008 2592 1008 0 FreeSans 480 90 0 0 I1/EN0
flabel metal3 2880 864 2880 864 0 FreeSans 480 90 0 0 I1/EN1
flabel metal3 4320 1008 4320 1008 0 FreeSans 480 90 0 0 I1/O
flabel metal2 2880 2016 2880 2016 0 FreeSans 960 0 0 0 I1/VSS
flabel metal2 2880 0 2880 0 0 FreeSans 960 0 0 0 I1/VDD
flabel space 1728 1008 1872 2016 0 FreeSans 320 90 0 0 I1/MN1_IBNDL0/nmos_boundary
flabel metal1 1266 1402 1326 1728 0 FreeSans 240 0 0 0 I1/MN0_IM0/S0
flabel metal1 1410 1402 1470 1728 0 FreeSans 240 0 0 0 I1/MN0_IM0/D0
flabel metal1 1554 1402 1614 1728 0 FreeSans 240 0 0 0 I1/MN0_IM0/S1
flabel metal1 1352 1260 1526 1332 0 FreeSans 240 0 0 0 I1/MN0_IM0/G0
rlabel pwell 1256 1340 1286 1362 5 I1/MN0_IM0/BODY
flabel space 1584 1008 1728 2016 0 FreeSans 320 90 0 0 I1/MN0_IBNDR0/nmos_boundary
flabel space 1152 1008 1296 2016 0 FreeSans 320 90 0 0 I1/MN0_IBNDL0/nmos_boundary
flabel space 1728 0 1872 1008 0 FreeSans 320 90 0 0 I1/MP1_IBNDL0/pmos_boundary
flabel metal1 1410 188 1470 594 0 FreeSans 160 0 0 0 I1/MP0_IM0/D0
flabel metal1 1352 684 1526 756 0 FreeSans 160 0 0 0 I1/MP0_IM0/G0
flabel metal1 1266 188 1326 594 0 FreeSans 160 0 0 0 I1/MP0_IM0/S0
flabel metal1 1554 188 1614 594 0 FreeSans 160 0 0 0 I1/MP0_IM0/S1
flabel nwell 1276 654 1300 670 0 FreeSans 80 0 0 0 I1/MP0_IM0/BODY
flabel space 1584 0 1728 1008 0 FreeSans 320 90 0 0 I1/MP0_IBNDR0/pmos_boundary
flabel space 1152 0 1296 1008 0 FreeSans 320 90 0 0 I1/MP0_IBNDL0/pmos_boundary
flabel space 2304 1008 2592 2016 0 FreeSans 320 90 0 0 I1/nspace0/NMOS_SPACE_2X
flabel metal1 1842 1402 1902 1728 0 FreeSans 240 0 0 0 I1/MN1_IM0/S0
flabel metal1 1986 1402 2046 1728 0 FreeSans 240 0 0 0 I1/MN1_IM0/D0
flabel metal1 2130 1402 2190 1728 0 FreeSans 240 0 0 0 I1/MN1_IM0/S1
flabel metal1 1928 1260 2102 1332 0 FreeSans 240 0 0 0 I1/MN1_IM0/G0
rlabel pwell 1832 1340 1862 1362 5 I1/MN1_IM0/BODY
flabel space 2160 1008 2304 2016 0 FreeSans 320 90 0 0 I1/MN1_IBNDR0/nmos_boundary
flabel space 2304 0 2592 1008 0 FreeSans 320 90 0 0 I1/pspace0/PMOS_SPACE_2X
flabel metal1 1986 188 2046 594 0 FreeSans 160 0 0 0 I1/MP1_IM0/D0
flabel metal1 1928 684 2102 756 0 FreeSans 160 0 0 0 I1/MP1_IM0/G0
flabel metal1 1842 188 1902 594 0 FreeSans 160 0 0 0 I1/MP1_IM0/S0
flabel metal1 2130 188 2190 594 0 FreeSans 160 0 0 0 I1/MP1_IM0/S1
flabel nwell 1852 654 1876 670 0 FreeSans 80 0 0 0 I1/MP1_IM0/BODY
flabel space 2160 0 2304 1008 0 FreeSans 320 90 0 0 I1/MP1_IBNDR0/pmos_boundary
flabel space 2592 1008 2880 2016 0 FreeSans 320 90 0 0 I1/nspace1/NMOS_SPACE_2X
flabel metal1 2994 1402 3054 1728 0 FreeSans 240 0 0 0 I1/MN2_IM0/S0
flabel metal1 3138 1402 3198 1728 0 FreeSans 240 0 0 0 I1/MN2_IM0/D0
flabel metal1 3282 1402 3342 1728 0 FreeSans 240 0 0 0 I1/MN2_IM0/S1
flabel metal1 3080 1260 3254 1332 0 FreeSans 240 0 0 0 I1/MN2_IM0/G0
rlabel pwell 2984 1340 3014 1362 5 I1/MN2_IM0/BODY
flabel space 2880 1008 3024 2016 0 FreeSans 320 90 0 0 I1/MN2_IBNDL0/nmos_boundary
flabel space 2592 0 2880 1008 0 FreeSans 320 90 0 0 I1/pspace1/PMOS_SPACE_2X
flabel metal1 3138 188 3198 594 0 FreeSans 160 0 0 0 I1/MP2_IM0/D0
flabel metal1 3080 684 3254 756 0 FreeSans 160 0 0 0 I1/MP2_IM0/G0
flabel metal1 2994 188 3054 594 0 FreeSans 160 0 0 0 I1/MP2_IM0/S0
flabel metal1 3282 188 3342 594 0 FreeSans 160 0 0 0 I1/MP2_IM0/S1
flabel nwell 3004 654 3028 670 0 FreeSans 80 0 0 0 I1/MP2_IM0/BODY
flabel space 2880 0 3024 1008 0 FreeSans 320 90 0 0 I1/MP2_IBNDL0/pmos_boundary
flabel metal1 3570 1402 3630 1728 0 FreeSans 240 0 0 0 I1/MN3_IM0/S0
flabel metal1 3714 1402 3774 1728 0 FreeSans 240 0 0 0 I1/MN3_IM0/D0
flabel metal1 3858 1402 3918 1728 0 FreeSans 240 0 0 0 I1/MN3_IM0/S1
flabel metal1 3656 1260 3830 1332 0 FreeSans 240 0 0 0 I1/MN3_IM0/G0
rlabel pwell 3560 1340 3590 1362 5 I1/MN3_IM0/BODY
flabel space 3456 1008 3600 2016 0 FreeSans 320 90 0 0 I1/MN3_IBNDL0/nmos_boundary
flabel space 3312 1008 3456 2016 0 FreeSans 320 90 0 0 I1/MN2_IBNDR0/nmos_boundary
flabel metal1 3714 188 3774 594 0 FreeSans 160 0 0 0 I1/MP3_IM0/D0
flabel metal1 3656 684 3830 756 0 FreeSans 160 0 0 0 I1/MP3_IM0/G0
flabel metal1 3570 188 3630 594 0 FreeSans 160 0 0 0 I1/MP3_IM0/S0
flabel metal1 3858 188 3918 594 0 FreeSans 160 0 0 0 I1/MP3_IM0/S1
flabel nwell 3580 654 3604 670 0 FreeSans 80 0 0 0 I1/MP3_IM0/BODY
flabel space 3456 0 3600 1008 0 FreeSans 320 90 0 0 I1/MP3_IBNDL0/pmos_boundary
flabel space 3312 0 3456 1008 0 FreeSans 320 90 0 0 I1/MP2_IBNDR0/pmos_boundary
flabel metal1 4146 1402 4206 1728 0 FreeSans 240 0 0 0 I1/MN4_IM0/S0
flabel metal1 4290 1402 4350 1728 0 FreeSans 240 0 0 0 I1/MN4_IM0/D0
flabel metal1 4434 1402 4494 1728 0 FreeSans 240 0 0 0 I1/MN4_IM0/S1
flabel metal1 4232 1260 4406 1332 0 FreeSans 240 0 0 0 I1/MN4_IM0/G0
rlabel pwell 4136 1340 4166 1362 5 I1/MN4_IM0/BODY
flabel space 4032 1008 4176 2016 0 FreeSans 320 90 0 0 I1/MN4_IBNDL0/nmos_boundary
flabel space 3888 1008 4032 2016 0 FreeSans 320 90 0 0 I1/MN3_IBNDR0/nmos_boundary
flabel metal1 4290 188 4350 594 0 FreeSans 160 0 0 0 I1/MP4_IM0/D0
flabel metal1 4232 684 4406 756 0 FreeSans 160 0 0 0 I1/MP4_IM0/G0
flabel metal1 4146 188 4206 594 0 FreeSans 160 0 0 0 I1/MP4_IM0/S0
flabel metal1 4434 188 4494 594 0 FreeSans 160 0 0 0 I1/MP4_IM0/S1
flabel nwell 4156 654 4180 670 0 FreeSans 80 0 0 0 I1/MP4_IM0/BODY
flabel space 4032 0 4176 1008 0 FreeSans 320 90 0 0 I1/MP4_IBNDL0/pmos_boundary
flabel space 3888 0 4032 1008 0 FreeSans 320 90 0 0 I1/MP3_IBNDR0/pmos_boundary
flabel space 4464 1008 4608 2016 0 FreeSans 320 90 0 0 I1/MN4_IBNDR0/nmos_boundary
flabel space 4464 0 4608 1008 0 FreeSans 320 90 0 0 I1/MP4_IBNDR0/pmos_boundary
flabel space 5040 0 5184 1024 0 FreeSans 320 90 0 0 I1/TAP0/MPT0_IBNDR0/ptap_boundary
flabel space 4608 0 4752 1024 0 FreeSans 320 90 0 0 I1/TAP0/MPT0_IBNDL0/ptap_boundary
flabel space 5040 992 5184 2016 0 FreeSans 320 90 0 0 I1/TAP0/MNT0_IBNDR0/ntap_boundary
flabel space 4608 992 4752 2016 0 FreeSans 320 90 0 0 I1/TAP0/MNT0_IBNDL0/ntap_boundary
flabel metal3 10800 3024 10800 3024 0 FreeSans 480 90 0 0 I3/I
flabel metal3 10944 3024 10944 3024 0 FreeSans 480 90 0 0 I3/O
flabel metal2 10944 2016 10944 2016 0 FreeSans 960 0 0 0 I3/VSS
flabel metal2 10944 4032 10944 4032 0 FreeSans 960 0 0 0 I3/VDD
flabel metal1 10914 3438 10974 3844 0 FreeSans 160 0 0 0 I3/MP0_IM0/D0
flabel metal1 10856 3276 11030 3348 0 FreeSans 160 0 0 0 I3/MP0_IM0/G0
flabel metal1 10770 3438 10830 3844 0 FreeSans 160 0 0 0 I3/MP0_IM0/S0
flabel metal1 11058 3438 11118 3844 0 FreeSans 160 0 0 0 I3/MP0_IM0/S1
flabel nwell 10780 3362 10804 3378 0 FreeSans 80 0 0 0 I3/MP0_IM0/BODY
flabel space 11088 3024 11232 4032 0 FreeSans 320 90 0 0 I3/MP0_IBNDR0/pmos_boundary
flabel space 10656 3024 10800 4032 0 FreeSans 320 90 0 0 I3/MP0_IBNDL0/pmos_boundary
flabel metal1 10770 2304 10830 2630 0 FreeSans 240 0 0 0 I3/MN0_IM0/S0
flabel metal1 10914 2304 10974 2630 0 FreeSans 240 0 0 0 I3/MN0_IM0/D0
flabel metal1 11058 2304 11118 2630 0 FreeSans 240 0 0 0 I3/MN0_IM0/S1
flabel metal1 10856 2700 11030 2772 0 FreeSans 240 0 0 0 I3/MN0_IM0/G0
rlabel pwell 10760 2670 10790 2692 1 I3/MN0_IM0/BODY
flabel space 11088 2016 11232 3024 0 FreeSans 320 90 0 0 I3/MN0_IBNDR0/nmos_boundary
flabel space 10656 2016 10800 3024 0 FreeSans 320 90 0 0 I3/MN0_IBNDL0/nmos_boundary
flabel space 11664 3008 11808 4032 0 FreeSans 320 90 0 0 TAP1_2/MPT0_IBNDR0/ptap_boundary
flabel space 11232 3008 11376 4032 0 FreeSans 320 90 0 0 TAP1_2/MPT0_IBNDL0/ptap_boundary
flabel space 11664 2016 11808 3040 0 FreeSans 320 90 0 0 TAP1_2/MNT0_IBNDR0/ntap_boundary
flabel space 11232 2016 11376 3040 0 FreeSans 320 90 0 0 TAP1_2/MNT0_IBNDL0/ntap_boundary
flabel metal3 12528 1008 12528 1008 0 FreeSans 480 90 0 0 I4/I
flabel metal3 12672 1008 12672 1008 0 FreeSans 480 90 0 0 I4/O
flabel metal2 12672 2016 12672 2016 0 FreeSans 960 0 0 0 I4/VSS
flabel metal2 12672 0 12672 0 0 FreeSans 960 0 0 0 I4/VDD
flabel metal1 12642 188 12702 594 0 FreeSans 160 0 0 0 I4/MP0_IM0/D0
flabel metal1 12584 684 12758 756 0 FreeSans 160 0 0 0 I4/MP0_IM0/G0
flabel metal1 12498 188 12558 594 0 FreeSans 160 0 0 0 I4/MP0_IM0/S0
flabel metal1 12786 188 12846 594 0 FreeSans 160 0 0 0 I4/MP0_IM0/S1
flabel nwell 12508 654 12532 670 0 FreeSans 80 0 0 0 I4/MP0_IM0/BODY
flabel space 12816 0 12960 1008 0 FreeSans 320 90 0 0 I4/MP0_IBNDR0/pmos_boundary
flabel space 12384 0 12528 1008 0 FreeSans 320 90 0 0 I4/MP0_IBNDL0/pmos_boundary
flabel metal1 12498 1402 12558 1728 0 FreeSans 240 0 0 0 I4/MN0_IM0/S0
flabel metal1 12642 1402 12702 1728 0 FreeSans 240 0 0 0 I4/MN0_IM0/D0
flabel metal1 12786 1402 12846 1728 0 FreeSans 240 0 0 0 I4/MN0_IM0/S1
flabel metal1 12584 1260 12758 1332 0 FreeSans 240 0 0 0 I4/MN0_IM0/G0
rlabel pwell 12488 1340 12518 1362 5 I4/MN0_IM0/BODY
flabel space 12816 1008 12960 2016 0 FreeSans 320 90 0 0 I4/MN0_IBNDR0/nmos_boundary
flabel space 12384 1008 12528 2016 0 FreeSans 320 90 0 0 I4/MN0_IBNDL0/nmos_boundary
flabel metal3 13104 1008 13104 1008 0 FreeSans 480 90 0 0 I5/I
flabel metal3 13248 1008 13248 1008 0 FreeSans 480 90 0 0 I5/O
flabel metal2 13248 2016 13248 2016 0 FreeSans 960 0 0 0 I5/VSS
flabel metal2 13248 0 13248 0 0 FreeSans 960 0 0 0 I5/VDD
flabel metal1 13218 188 13278 594 0 FreeSans 160 0 0 0 I5/MP0_IM0/D0
flabel metal1 13160 684 13334 756 0 FreeSans 160 0 0 0 I5/MP0_IM0/G0
flabel metal1 13074 188 13134 594 0 FreeSans 160 0 0 0 I5/MP0_IM0/S0
flabel metal1 13362 188 13422 594 0 FreeSans 160 0 0 0 I5/MP0_IM0/S1
flabel nwell 13084 654 13108 670 0 FreeSans 80 0 0 0 I5/MP0_IM0/BODY
flabel space 13392 0 13536 1008 0 FreeSans 320 90 0 0 I5/MP0_IBNDR0/pmos_boundary
flabel space 12960 0 13104 1008 0 FreeSans 320 90 0 0 I5/MP0_IBNDL0/pmos_boundary
flabel metal1 13074 1402 13134 1728 0 FreeSans 240 0 0 0 I5/MN0_IM0/S0
flabel metal1 13218 1402 13278 1728 0 FreeSans 240 0 0 0 I5/MN0_IM0/D0
flabel metal1 13362 1402 13422 1728 0 FreeSans 240 0 0 0 I5/MN0_IM0/S1
flabel metal1 13160 1260 13334 1332 0 FreeSans 240 0 0 0 I5/MN0_IM0/G0
rlabel pwell 13064 1340 13094 1362 5 I5/MN0_IM0/BODY
flabel space 13392 1008 13536 2016 0 FreeSans 320 90 0 0 I5/MN0_IBNDR0/nmos_boundary
flabel space 12960 1008 13104 2016 0 FreeSans 320 90 0 0 I5/MN0_IBNDL0/nmos_boundary
flabel metal3 12096 3024 12096 3024 0 FreeSans 480 90 0 0 I21/I0
flabel metal3 14400 3024 14400 3024 0 FreeSans 480 90 0 0 I21/I1
flabel metal3 13248 3024 13248 3024 0 FreeSans 480 90 0 0 I21/EN0
flabel metal3 13536 3168 13536 3168 0 FreeSans 480 90 0 0 I21/EN1
flabel metal3 14976 3024 14976 3024 0 FreeSans 480 90 0 0 I21/O
flabel metal2 13536 2016 13536 2016 0 FreeSans 960 0 0 0 I21/VSS
flabel metal2 13536 4032 13536 4032 0 FreeSans 960 0 0 0 I21/VDD
flabel space 12384 2016 12528 3024 0 FreeSans 320 90 0 0 I21/MN1_IBNDL0/nmos_boundary
flabel metal1 11922 2304 11982 2630 0 FreeSans 240 0 0 0 I21/MN0_IM0/S0
flabel metal1 12066 2304 12126 2630 0 FreeSans 240 0 0 0 I21/MN0_IM0/D0
flabel metal1 12210 2304 12270 2630 0 FreeSans 240 0 0 0 I21/MN0_IM0/S1
flabel metal1 12008 2700 12182 2772 0 FreeSans 240 0 0 0 I21/MN0_IM0/G0
rlabel pwell 11912 2670 11942 2692 1 I21/MN0_IM0/BODY
flabel space 12240 2016 12384 3024 0 FreeSans 320 90 0 0 I21/MN0_IBNDR0/nmos_boundary
flabel space 11808 2016 11952 3024 0 FreeSans 320 90 0 0 I21/MN0_IBNDL0/nmos_boundary
flabel space 12384 3024 12528 4032 0 FreeSans 320 90 0 0 I21/MP1_IBNDL0/pmos_boundary
flabel metal1 12066 3438 12126 3844 0 FreeSans 160 0 0 0 I21/MP0_IM0/D0
flabel metal1 12008 3276 12182 3348 0 FreeSans 160 0 0 0 I21/MP0_IM0/G0
flabel metal1 11922 3438 11982 3844 0 FreeSans 160 0 0 0 I21/MP0_IM0/S0
flabel metal1 12210 3438 12270 3844 0 FreeSans 160 0 0 0 I21/MP0_IM0/S1
flabel nwell 11932 3362 11956 3378 0 FreeSans 80 0 0 0 I21/MP0_IM0/BODY
flabel space 12240 3024 12384 4032 0 FreeSans 320 90 0 0 I21/MP0_IBNDR0/pmos_boundary
flabel space 11808 3024 11952 4032 0 FreeSans 320 90 0 0 I21/MP0_IBNDL0/pmos_boundary
flabel space 12960 2016 13248 3024 0 FreeSans 320 90 0 0 I21/nspace0/NMOS_SPACE_2X
flabel metal1 12498 2304 12558 2630 0 FreeSans 240 0 0 0 I21/MN1_IM0/S0
flabel metal1 12642 2304 12702 2630 0 FreeSans 240 0 0 0 I21/MN1_IM0/D0
flabel metal1 12786 2304 12846 2630 0 FreeSans 240 0 0 0 I21/MN1_IM0/S1
flabel metal1 12584 2700 12758 2772 0 FreeSans 240 0 0 0 I21/MN1_IM0/G0
rlabel pwell 12488 2670 12518 2692 1 I21/MN1_IM0/BODY
flabel space 12816 2016 12960 3024 0 FreeSans 320 90 0 0 I21/MN1_IBNDR0/nmos_boundary
flabel space 12960 3024 13248 4032 0 FreeSans 320 90 0 0 I21/pspace0/PMOS_SPACE_2X
flabel metal1 12642 3438 12702 3844 0 FreeSans 160 0 0 0 I21/MP1_IM0/D0
flabel metal1 12584 3276 12758 3348 0 FreeSans 160 0 0 0 I21/MP1_IM0/G0
flabel metal1 12498 3438 12558 3844 0 FreeSans 160 0 0 0 I21/MP1_IM0/S0
flabel metal1 12786 3438 12846 3844 0 FreeSans 160 0 0 0 I21/MP1_IM0/S1
flabel nwell 12508 3362 12532 3378 0 FreeSans 80 0 0 0 I21/MP1_IM0/BODY
flabel space 12816 3024 12960 4032 0 FreeSans 320 90 0 0 I21/MP1_IBNDR0/pmos_boundary
flabel space 13248 2016 13536 3024 0 FreeSans 320 90 0 0 I21/nspace1/NMOS_SPACE_2X
flabel metal1 13650 2304 13710 2630 0 FreeSans 240 0 0 0 I21/MN2_IM0/S0
flabel metal1 13794 2304 13854 2630 0 FreeSans 240 0 0 0 I21/MN2_IM0/D0
flabel metal1 13938 2304 13998 2630 0 FreeSans 240 0 0 0 I21/MN2_IM0/S1
flabel metal1 13736 2700 13910 2772 0 FreeSans 240 0 0 0 I21/MN2_IM0/G0
rlabel pwell 13640 2670 13670 2692 1 I21/MN2_IM0/BODY
flabel space 13536 2016 13680 3024 0 FreeSans 320 90 0 0 I21/MN2_IBNDL0/nmos_boundary
flabel space 13248 3024 13536 4032 0 FreeSans 320 90 0 0 I21/pspace1/PMOS_SPACE_2X
flabel metal1 13794 3438 13854 3844 0 FreeSans 160 0 0 0 I21/MP2_IM0/D0
flabel metal1 13736 3276 13910 3348 0 FreeSans 160 0 0 0 I21/MP2_IM0/G0
flabel metal1 13650 3438 13710 3844 0 FreeSans 160 0 0 0 I21/MP2_IM0/S0
flabel metal1 13938 3438 13998 3844 0 FreeSans 160 0 0 0 I21/MP2_IM0/S1
flabel nwell 13660 3362 13684 3378 0 FreeSans 80 0 0 0 I21/MP2_IM0/BODY
flabel space 13536 3024 13680 4032 0 FreeSans 320 90 0 0 I21/MP2_IBNDL0/pmos_boundary
flabel metal1 14226 2304 14286 2630 0 FreeSans 240 0 0 0 I21/MN3_IM0/S0
flabel metal1 14370 2304 14430 2630 0 FreeSans 240 0 0 0 I21/MN3_IM0/D0
flabel metal1 14514 2304 14574 2630 0 FreeSans 240 0 0 0 I21/MN3_IM0/S1
flabel metal1 14312 2700 14486 2772 0 FreeSans 240 0 0 0 I21/MN3_IM0/G0
rlabel pwell 14216 2670 14246 2692 1 I21/MN3_IM0/BODY
flabel space 14112 2016 14256 3024 0 FreeSans 320 90 0 0 I21/MN3_IBNDL0/nmos_boundary
flabel space 13968 2016 14112 3024 0 FreeSans 320 90 0 0 I21/MN2_IBNDR0/nmos_boundary
flabel metal1 14370 3438 14430 3844 0 FreeSans 160 0 0 0 I21/MP3_IM0/D0
flabel metal1 14312 3276 14486 3348 0 FreeSans 160 0 0 0 I21/MP3_IM0/G0
flabel metal1 14226 3438 14286 3844 0 FreeSans 160 0 0 0 I21/MP3_IM0/S0
flabel metal1 14514 3438 14574 3844 0 FreeSans 160 0 0 0 I21/MP3_IM0/S1
flabel nwell 14236 3362 14260 3378 0 FreeSans 80 0 0 0 I21/MP3_IM0/BODY
flabel space 14112 3024 14256 4032 0 FreeSans 320 90 0 0 I21/MP3_IBNDL0/pmos_boundary
flabel space 13968 3024 14112 4032 0 FreeSans 320 90 0 0 I21/MP2_IBNDR0/pmos_boundary
flabel metal1 14802 2304 14862 2630 0 FreeSans 240 0 0 0 I21/MN4_IM0/S0
flabel metal1 14946 2304 15006 2630 0 FreeSans 240 0 0 0 I21/MN4_IM0/D0
flabel metal1 15090 2304 15150 2630 0 FreeSans 240 0 0 0 I21/MN4_IM0/S1
flabel metal1 14888 2700 15062 2772 0 FreeSans 240 0 0 0 I21/MN4_IM0/G0
rlabel pwell 14792 2670 14822 2692 1 I21/MN4_IM0/BODY
flabel space 14688 2016 14832 3024 0 FreeSans 320 90 0 0 I21/MN4_IBNDL0/nmos_boundary
flabel space 14544 2016 14688 3024 0 FreeSans 320 90 0 0 I21/MN3_IBNDR0/nmos_boundary
flabel metal1 14946 3438 15006 3844 0 FreeSans 160 0 0 0 I21/MP4_IM0/D0
flabel metal1 14888 3276 15062 3348 0 FreeSans 160 0 0 0 I21/MP4_IM0/G0
flabel metal1 14802 3438 14862 3844 0 FreeSans 160 0 0 0 I21/MP4_IM0/S0
flabel metal1 15090 3438 15150 3844 0 FreeSans 160 0 0 0 I21/MP4_IM0/S1
flabel nwell 14812 3362 14836 3378 0 FreeSans 80 0 0 0 I21/MP4_IM0/BODY
flabel space 14688 3024 14832 4032 0 FreeSans 320 90 0 0 I21/MP4_IBNDL0/pmos_boundary
flabel space 14544 3024 14688 4032 0 FreeSans 320 90 0 0 I21/MP3_IBNDR0/pmos_boundary
flabel space 15120 2016 15264 3024 0 FreeSans 320 90 0 0 I21/MN4_IBNDR0/nmos_boundary
flabel space 15120 3024 15264 4032 0 FreeSans 320 90 0 0 I21/MP4_IBNDR0/pmos_boundary
flabel space 15696 3008 15840 4032 0 FreeSans 320 90 0 0 I21/TAP0/MPT0_IBNDR0/ptap_boundary
flabel space 15264 3008 15408 4032 0 FreeSans 320 90 0 0 I21/TAP0/MPT0_IBNDL0/ptap_boundary
flabel space 15696 2016 15840 3040 0 FreeSans 320 90 0 0 I21/TAP0/MNT0_IBNDR0/ntap_boundary
flabel space 15264 2016 15408 3040 0 FreeSans 320 90 0 0 I21/TAP0/MNT0_IBNDL0/ntap_boundary
flabel metal3 13680 1008 13680 1008 0 FreeSans 480 90 0 0 I6/I
flabel metal3 13824 1008 13824 1008 0 FreeSans 480 90 0 0 I6/O
flabel metal2 13824 2016 13824 2016 0 FreeSans 960 0 0 0 I6/VSS
flabel metal2 13824 0 13824 0 0 FreeSans 960 0 0 0 I6/VDD
flabel metal1 13794 188 13854 594 0 FreeSans 160 0 0 0 I6/MP0_IM0/D0
flabel metal1 13736 684 13910 756 0 FreeSans 160 0 0 0 I6/MP0_IM0/G0
flabel metal1 13650 188 13710 594 0 FreeSans 160 0 0 0 I6/MP0_IM0/S0
flabel metal1 13938 188 13998 594 0 FreeSans 160 0 0 0 I6/MP0_IM0/S1
flabel nwell 13660 654 13684 670 0 FreeSans 80 0 0 0 I6/MP0_IM0/BODY
flabel space 13968 0 14112 1008 0 FreeSans 320 90 0 0 I6/MP0_IBNDR0/pmos_boundary
flabel space 13536 0 13680 1008 0 FreeSans 320 90 0 0 I6/MP0_IBNDL0/pmos_boundary
flabel metal1 13650 1402 13710 1728 0 FreeSans 240 0 0 0 I6/MN0_IM0/S0
flabel metal1 13794 1402 13854 1728 0 FreeSans 240 0 0 0 I6/MN0_IM0/D0
flabel metal1 13938 1402 13998 1728 0 FreeSans 240 0 0 0 I6/MN0_IM0/S1
flabel metal1 13736 1260 13910 1332 0 FreeSans 240 0 0 0 I6/MN0_IM0/G0
rlabel pwell 13640 1340 13670 1362 5 I6/MN0_IM0/BODY
flabel space 13968 1008 14112 2016 0 FreeSans 320 90 0 0 I6/MN0_IBNDR0/nmos_boundary
flabel space 13536 1008 13680 2016 0 FreeSans 320 90 0 0 I6/MN0_IBNDL0/nmos_boundary
flabel space 14544 0 14688 1024 0 FreeSans 320 90 0 0 TAP0_2/MPT0_IBNDR0/ptap_boundary
flabel space 14112 0 14256 1024 0 FreeSans 320 90 0 0 TAP0_2/MPT0_IBNDL0/ptap_boundary
flabel space 14544 992 14688 2016 0 FreeSans 320 90 0 0 TAP0_2/MNT0_IBNDR0/ntap_boundary
flabel space 14112 992 14256 2016 0 FreeSans 320 90 0 0 TAP0_2/MNT0_IBNDL0/ntap_boundary
flabel metal3 14832 1008 14832 1008 0 FreeSans 480 90 0 0 I7/I
flabel metal3 14976 1008 14976 1008 0 FreeSans 480 90 0 0 I7/O
flabel metal2 14976 2016 14976 2016 0 FreeSans 960 0 0 0 I7/VSS
flabel metal2 14976 0 14976 0 0 FreeSans 960 0 0 0 I7/VDD
flabel metal1 14946 188 15006 594 0 FreeSans 160 0 0 0 I7/MP0_IM0/D0
flabel metal1 14888 684 15062 756 0 FreeSans 160 0 0 0 I7/MP0_IM0/G0
flabel metal1 14802 188 14862 594 0 FreeSans 160 0 0 0 I7/MP0_IM0/S0
flabel metal1 15090 188 15150 594 0 FreeSans 160 0 0 0 I7/MP0_IM0/S1
flabel nwell 14812 654 14836 670 0 FreeSans 80 0 0 0 I7/MP0_IM0/BODY
flabel space 15120 0 15264 1008 0 FreeSans 320 90 0 0 I7/MP0_IBNDR0/pmos_boundary
flabel space 14688 0 14832 1008 0 FreeSans 320 90 0 0 I7/MP0_IBNDL0/pmos_boundary
flabel metal1 14802 1402 14862 1728 0 FreeSans 240 0 0 0 I7/MN0_IM0/S0
flabel metal1 14946 1402 15006 1728 0 FreeSans 240 0 0 0 I7/MN0_IM0/D0
flabel metal1 15090 1402 15150 1728 0 FreeSans 240 0 0 0 I7/MN0_IM0/S1
flabel metal1 14888 1260 15062 1332 0 FreeSans 240 0 0 0 I7/MN0_IM0/G0
rlabel pwell 14792 1340 14822 1362 5 I7/MN0_IM0/BODY
flabel space 15120 1008 15264 2016 0 FreeSans 320 90 0 0 I7/MN0_IBNDR0/nmos_boundary
flabel space 14688 1008 14832 2016 0 FreeSans 320 90 0 0 I7/MN0_IBNDL0/nmos_boundary
flabel metal3 15696 1008 15696 1008 0 FreeSans 480 90 0 0 I22/I
flabel metal3 15552 1008 15552 1008 0 FreeSans 480 90 0 0 I22/O
flabel metal2 15552 2016 15552 2016 0 FreeSans 960 0 0 0 I22/VSS
flabel metal2 15552 0 15552 0 0 FreeSans 960 0 0 0 I22/VDD
flabel metal1 15522 188 15582 594 0 FreeSans 160 0 0 0 I22/MP0_IM0/D0
flabel metal1 15466 684 15640 756 0 FreeSans 160 0 0 0 I22/MP0_IM0/G0
flabel metal1 15666 188 15726 594 0 FreeSans 160 0 0 0 I22/MP0_IM0/S0
flabel metal1 15378 188 15438 594 0 FreeSans 160 0 0 0 I22/MP0_IM0/S1
flabel nwell 15692 654 15716 670 0 FreeSans 80 0 0 0 I22/MP0_IM0/BODY
flabel space 15264 0 15408 1008 0 FreeSans 320 90 0 0 I22/MP0_IBNDR0/pmos_boundary
flabel space 15696 0 15840 1008 0 FreeSans 320 90 0 0 I22/MP0_IBNDL0/pmos_boundary
flabel metal1 15666 1402 15726 1728 0 FreeSans 240 0 0 0 I22/MN0_IM0/S0
flabel metal1 15522 1402 15582 1728 0 FreeSans 240 0 0 0 I22/MN0_IM0/D0
flabel metal1 15378 1402 15438 1728 0 FreeSans 240 0 0 0 I22/MN0_IM0/S1
flabel metal1 15466 1260 15640 1332 0 FreeSans 240 0 0 0 I22/MN0_IM0/G0
rlabel pwell 15706 1340 15736 1362 5 I22/MN0_IM0/BODY
flabel space 15264 1008 15408 2016 0 FreeSans 320 90 0 0 I22/MN0_IBNDR0/nmos_boundary
flabel space 15696 1008 15840 2016 0 FreeSans 320 90 0 0 I22/MN0_IBNDL0/nmos_boundary
flabel metal3 15984 1008 15984 1008 0 FreeSans 480 90 0 0 I23/I
flabel metal3 16416 1008 16416 1008 0 FreeSans 480 90 0 0 I23/O
flabel metal2 16272 2016 16272 2016 0 FreeSans 960 0 0 0 I23/VSS
flabel metal2 16272 0 16272 0 0 FreeSans 960 0 0 0 I23/VDD
flabel metal1 16098 188 16158 594 0 FreeSans 160 0 0 0 I23/MP0_IM0[0]/D0
flabel metal1 16040 684 16214 756 0 FreeSans 160 0 0 0 I23/MP0_IM0[0]/G0
flabel metal1 15954 188 16014 594 0 FreeSans 160 0 0 0 I23/MP0_IM0[0]/S0
flabel metal1 16242 188 16302 594 0 FreeSans 160 0 0 0 I23/MP0_IM0[0]/S1
flabel nwell 15964 654 15988 670 0 FreeSans 80 0 0 0 I23/MP0_IM0[0]/BODY
flabel metal1 16386 188 16446 594 0 FreeSans 160 0 0 0 I23/MP0_IM0[1]/D0
flabel metal1 16328 684 16502 756 0 FreeSans 160 0 0 0 I23/MP0_IM0[1]/G0
flabel metal1 16242 188 16302 594 0 FreeSans 160 0 0 0 I23/MP0_IM0[1]/S0
flabel metal1 16530 188 16590 594 0 FreeSans 160 0 0 0 I23/MP0_IM0[1]/S1
flabel nwell 16252 654 16276 670 0 FreeSans 80 0 0 0 I23/MP0_IM0[1]/BODY
flabel space 16560 0 16704 1008 0 FreeSans 320 90 0 0 I23/MP0_IBNDR0/pmos_boundary
flabel space 15840 0 15984 1008 0 FreeSans 320 90 0 0 I23/MP0_IBNDL0/pmos_boundary
flabel metal1 15954 1402 16014 1728 0 FreeSans 240 0 0 0 I23/MN0_IM0[0]/S0
flabel metal1 16098 1402 16158 1728 0 FreeSans 240 0 0 0 I23/MN0_IM0[0]/D0
flabel metal1 16242 1402 16302 1728 0 FreeSans 240 0 0 0 I23/MN0_IM0[0]/S1
flabel metal1 16040 1260 16214 1332 0 FreeSans 240 0 0 0 I23/MN0_IM0[0]/G0
rlabel pwell 15944 1340 15974 1362 5 I23/MN0_IM0[0]/BODY
flabel metal1 16242 1402 16302 1728 0 FreeSans 240 0 0 0 I23/MN0_IM0[1]/S0
flabel metal1 16386 1402 16446 1728 0 FreeSans 240 0 0 0 I23/MN0_IM0[1]/D0
flabel metal1 16530 1402 16590 1728 0 FreeSans 240 0 0 0 I23/MN0_IM0[1]/S1
flabel metal1 16328 1260 16502 1332 0 FreeSans 240 0 0 0 I23/MN0_IM0[1]/G0
rlabel pwell 16232 1340 16262 1362 5 I23/MN0_IM0[1]/BODY
flabel space 16560 1008 16704 2016 0 FreeSans 320 90 0 0 I23/MN0_IBNDR0/nmos_boundary
flabel space 15840 1008 15984 2016 0 FreeSans 320 90 0 0 I23/MN0_IBNDL0/nmos_boundary
flabel space 16272 3008 16416 4032 0 FreeSans 320 90 0 0 TAP1_3/MPT0_IBNDR0/ptap_boundary
flabel space 15840 3008 15984 4032 0 FreeSans 320 90 0 0 TAP1_3/MPT0_IBNDL0/ptap_boundary
flabel space 16272 2016 16416 3040 0 FreeSans 320 90 0 0 TAP1_3/MNT0_IBNDR0/ntap_boundary
flabel space 15840 2016 15984 3040 0 FreeSans 320 90 0 0 TAP1_3/MNT0_IBNDL0/ntap_boundary
flabel space 17136 0 17280 1024 0 FreeSans 320 90 0 0 TAP0_3/MPT0_IBNDR0/ptap_boundary
flabel space 16704 0 16848 1024 0 FreeSans 320 90 0 0 TAP0_3/MPT0_IBNDL0/ptap_boundary
flabel space 17136 992 17280 2016 0 FreeSans 320 90 0 0 TAP0_3/MNT0_IBNDR0/ntap_boundary
flabel space 16704 992 16848 2016 0 FreeSans 320 90 0 0 TAP0_3/MNT0_IBNDL0/ntap_boundary
flabel metal3 17424 1008 17424 1008 0 FreeSans 480 90 0 0 I24/I
flabel metal3 20736 1008 20736 1008 0 FreeSans 480 90 0 0 I24/O
flabel metal2 19152 2016 19152 2016 0 FreeSans 960 0 0 0 I24/VSS
flabel metal2 19152 0 19152 0 0 FreeSans 960 0 0 0 I24/VDD
flabel metal1 17538 188 17598 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[0]/D0
flabel metal1 17480 684 17654 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[0]/G0
flabel metal1 17394 188 17454 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[0]/S0
flabel metal1 17682 188 17742 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[0]/S1
flabel nwell 17404 654 17428 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[0]/BODY
flabel metal1 17826 188 17886 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[1]/D0
flabel metal1 17768 684 17942 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[1]/G0
flabel metal1 17682 188 17742 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[1]/S0
flabel metal1 17970 188 18030 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[1]/S1
flabel nwell 17692 654 17716 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[1]/BODY
flabel metal1 18114 188 18174 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[2]/D0
flabel metal1 18056 684 18230 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[2]/G0
flabel metal1 17970 188 18030 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[2]/S0
flabel metal1 18258 188 18318 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[2]/S1
flabel nwell 17980 654 18004 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[2]/BODY
flabel metal1 18402 188 18462 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[3]/D0
flabel metal1 18344 684 18518 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[3]/G0
flabel metal1 18258 188 18318 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[3]/S0
flabel metal1 18546 188 18606 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[3]/S1
flabel nwell 18268 654 18292 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[3]/BODY
flabel metal1 18690 188 18750 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[4]/D0
flabel metal1 18632 684 18806 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[4]/G0
flabel metal1 18546 188 18606 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[4]/S0
flabel metal1 18834 188 18894 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[4]/S1
flabel nwell 18556 654 18580 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[4]/BODY
flabel metal1 18978 188 19038 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[5]/D0
flabel metal1 18920 684 19094 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[5]/G0
flabel metal1 18834 188 18894 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[5]/S0
flabel metal1 19122 188 19182 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[5]/S1
flabel nwell 18844 654 18868 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[5]/BODY
flabel metal1 19266 188 19326 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[6]/D0
flabel metal1 19208 684 19382 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[6]/G0
flabel metal1 19122 188 19182 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[6]/S0
flabel metal1 19410 188 19470 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[6]/S1
flabel nwell 19132 654 19156 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[6]/BODY
flabel metal1 19554 188 19614 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[7]/D0
flabel metal1 19496 684 19670 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[7]/G0
flabel metal1 19410 188 19470 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[7]/S0
flabel metal1 19698 188 19758 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[7]/S1
flabel nwell 19420 654 19444 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[7]/BODY
flabel metal1 19842 188 19902 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[8]/D0
flabel metal1 19784 684 19958 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[8]/G0
flabel metal1 19698 188 19758 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[8]/S0
flabel metal1 19986 188 20046 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[8]/S1
flabel nwell 19708 654 19732 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[8]/BODY
flabel metal1 20130 188 20190 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[9]/D0
flabel metal1 20072 684 20246 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[9]/G0
flabel metal1 19986 188 20046 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[9]/S0
flabel metal1 20274 188 20334 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[9]/S1
flabel nwell 19996 654 20020 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[9]/BODY
flabel metal1 20418 188 20478 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[10]/D0
flabel metal1 20360 684 20534 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[10]/G0
flabel metal1 20274 188 20334 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[10]/S0
flabel metal1 20562 188 20622 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[10]/S1
flabel nwell 20284 654 20308 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[10]/BODY
flabel metal1 20706 188 20766 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[11]/D0
flabel metal1 20648 684 20822 756 0 FreeSans 160 0 0 0 I24/MP0_IM0[11]/G0
flabel metal1 20562 188 20622 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[11]/S0
flabel metal1 20850 188 20910 594 0 FreeSans 160 0 0 0 I24/MP0_IM0[11]/S1
flabel nwell 20572 654 20596 670 0 FreeSans 80 0 0 0 I24/MP0_IM0[11]/BODY
flabel space 20880 0 21024 1008 0 FreeSans 320 90 0 0 I24/MP0_IBNDR0/pmos_boundary
flabel space 17280 0 17424 1008 0 FreeSans 320 90 0 0 I24/MP0_IBNDL0/pmos_boundary
flabel metal1 17394 1402 17454 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[0]/S0
flabel metal1 17538 1402 17598 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[0]/D0
flabel metal1 17682 1402 17742 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[0]/S1
flabel metal1 17480 1260 17654 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[0]/G0
rlabel pwell 17384 1340 17414 1362 5 I24/MN0_IM0[0]/BODY
flabel metal1 17682 1402 17742 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[1]/S0
flabel metal1 17826 1402 17886 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[1]/D0
flabel metal1 17970 1402 18030 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[1]/S1
flabel metal1 17768 1260 17942 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[1]/G0
rlabel pwell 17672 1340 17702 1362 5 I24/MN0_IM0[1]/BODY
flabel metal1 17970 1402 18030 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[2]/S0
flabel metal1 18114 1402 18174 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[2]/D0
flabel metal1 18258 1402 18318 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[2]/S1
flabel metal1 18056 1260 18230 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[2]/G0
rlabel pwell 17960 1340 17990 1362 5 I24/MN0_IM0[2]/BODY
flabel metal1 18258 1402 18318 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[3]/S0
flabel metal1 18402 1402 18462 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[3]/D0
flabel metal1 18546 1402 18606 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[3]/S1
flabel metal1 18344 1260 18518 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[3]/G0
rlabel pwell 18248 1340 18278 1362 5 I24/MN0_IM0[3]/BODY
flabel metal1 18546 1402 18606 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[4]/S0
flabel metal1 18690 1402 18750 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[4]/D0
flabel metal1 18834 1402 18894 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[4]/S1
flabel metal1 18632 1260 18806 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[4]/G0
rlabel pwell 18536 1340 18566 1362 5 I24/MN0_IM0[4]/BODY
flabel metal1 18834 1402 18894 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[5]/S0
flabel metal1 18978 1402 19038 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[5]/D0
flabel metal1 19122 1402 19182 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[5]/S1
flabel metal1 18920 1260 19094 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[5]/G0
rlabel pwell 18824 1340 18854 1362 5 I24/MN0_IM0[5]/BODY
flabel metal1 19122 1402 19182 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[6]/S0
flabel metal1 19266 1402 19326 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[6]/D0
flabel metal1 19410 1402 19470 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[6]/S1
flabel metal1 19208 1260 19382 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[6]/G0
rlabel pwell 19112 1340 19142 1362 5 I24/MN0_IM0[6]/BODY
flabel metal1 19410 1402 19470 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[7]/S0
flabel metal1 19554 1402 19614 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[7]/D0
flabel metal1 19698 1402 19758 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[7]/S1
flabel metal1 19496 1260 19670 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[7]/G0
rlabel pwell 19400 1340 19430 1362 5 I24/MN0_IM0[7]/BODY
flabel metal1 19698 1402 19758 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[8]/S0
flabel metal1 19842 1402 19902 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[8]/D0
flabel metal1 19986 1402 20046 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[8]/S1
flabel metal1 19784 1260 19958 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[8]/G0
rlabel pwell 19688 1340 19718 1362 5 I24/MN0_IM0[8]/BODY
flabel metal1 19986 1402 20046 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[9]/S0
flabel metal1 20130 1402 20190 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[9]/D0
flabel metal1 20274 1402 20334 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[9]/S1
flabel metal1 20072 1260 20246 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[9]/G0
rlabel pwell 19976 1340 20006 1362 5 I24/MN0_IM0[9]/BODY
flabel metal1 20274 1402 20334 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[10]/S0
flabel metal1 20418 1402 20478 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[10]/D0
flabel metal1 20562 1402 20622 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[10]/S1
flabel metal1 20360 1260 20534 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[10]/G0
rlabel pwell 20264 1340 20294 1362 5 I24/MN0_IM0[10]/BODY
flabel metal1 20562 1402 20622 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[11]/S0
flabel metal1 20706 1402 20766 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[11]/D0
flabel metal1 20850 1402 20910 1728 0 FreeSans 240 0 0 0 I24/MN0_IM0[11]/S1
flabel metal1 20648 1260 20822 1332 0 FreeSans 240 0 0 0 I24/MN0_IM0[11]/G0
rlabel pwell 20552 1340 20582 1362 5 I24/MN0_IM0[11]/BODY
flabel space 20880 1008 21024 2016 0 FreeSans 320 90 0 0 I24/MN0_IBNDR0/nmos_boundary
flabel space 17280 1008 17424 2016 0 FreeSans 320 90 0 0 I24/MN0_IBNDL0/nmos_boundary
flabel metal3 20016 3024 20016 3024 0 FreeSans 480 90 0 0 I14/I
flabel metal3 16704 3024 16704 3024 0 FreeSans 480 90 0 0 I14/O
flabel metal2 18288 2016 18288 2016 0 FreeSans 960 0 0 0 I14/VSS
flabel metal2 18288 4032 18288 4032 0 FreeSans 960 0 0 0 I14/VDD
flabel metal1 19842 3438 19902 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[0]/D0
flabel metal1 19786 3276 19960 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[0]/G0
flabel metal1 19986 3438 20046 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[0]/S0
flabel metal1 19698 3438 19758 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[0]/S1
flabel nwell 20012 3362 20036 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[0]/BODY
flabel metal1 19554 3438 19614 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[1]/D0
flabel metal1 19498 3276 19672 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[1]/G0
flabel metal1 19698 3438 19758 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[1]/S0
flabel metal1 19410 3438 19470 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[1]/S1
flabel nwell 19724 3362 19748 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[1]/BODY
flabel metal1 19266 3438 19326 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[2]/D0
flabel metal1 19210 3276 19384 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[2]/G0
flabel metal1 19410 3438 19470 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[2]/S0
flabel metal1 19122 3438 19182 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[2]/S1
flabel nwell 19436 3362 19460 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[2]/BODY
flabel metal1 18978 3438 19038 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[3]/D0
flabel metal1 18922 3276 19096 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[3]/G0
flabel metal1 19122 3438 19182 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[3]/S0
flabel metal1 18834 3438 18894 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[3]/S1
flabel nwell 19148 3362 19172 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[3]/BODY
flabel metal1 18690 3438 18750 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[4]/D0
flabel metal1 18634 3276 18808 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[4]/G0
flabel metal1 18834 3438 18894 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[4]/S0
flabel metal1 18546 3438 18606 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[4]/S1
flabel nwell 18860 3362 18884 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[4]/BODY
flabel metal1 18402 3438 18462 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[5]/D0
flabel metal1 18346 3276 18520 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[5]/G0
flabel metal1 18546 3438 18606 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[5]/S0
flabel metal1 18258 3438 18318 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[5]/S1
flabel nwell 18572 3362 18596 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[5]/BODY
flabel metal1 18114 3438 18174 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[6]/D0
flabel metal1 18058 3276 18232 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[6]/G0
flabel metal1 18258 3438 18318 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[6]/S0
flabel metal1 17970 3438 18030 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[6]/S1
flabel nwell 18284 3362 18308 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[6]/BODY
flabel metal1 17826 3438 17886 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[7]/D0
flabel metal1 17770 3276 17944 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[7]/G0
flabel metal1 17970 3438 18030 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[7]/S0
flabel metal1 17682 3438 17742 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[7]/S1
flabel nwell 17996 3362 18020 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[7]/BODY
flabel metal1 17538 3438 17598 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[8]/D0
flabel metal1 17482 3276 17656 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[8]/G0
flabel metal1 17682 3438 17742 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[8]/S0
flabel metal1 17394 3438 17454 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[8]/S1
flabel nwell 17708 3362 17732 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[8]/BODY
flabel metal1 17250 3438 17310 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[9]/D0
flabel metal1 17194 3276 17368 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[9]/G0
flabel metal1 17394 3438 17454 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[9]/S0
flabel metal1 17106 3438 17166 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[9]/S1
flabel nwell 17420 3362 17444 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[9]/BODY
flabel metal1 16962 3438 17022 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[10]/D0
flabel metal1 16906 3276 17080 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[10]/G0
flabel metal1 17106 3438 17166 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[10]/S0
flabel metal1 16818 3438 16878 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[10]/S1
flabel nwell 17132 3362 17156 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[10]/BODY
flabel metal1 16674 3438 16734 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[11]/D0
flabel metal1 16618 3276 16792 3348 0 FreeSans 160 0 0 0 I14/MP0_IM0[11]/G0
flabel metal1 16818 3438 16878 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[11]/S0
flabel metal1 16530 3438 16590 3844 0 FreeSans 160 0 0 0 I14/MP0_IM0[11]/S1
flabel nwell 16844 3362 16868 3378 0 FreeSans 80 0 0 0 I14/MP0_IM0[11]/BODY
flabel space 16416 3024 16560 4032 0 FreeSans 320 90 0 0 I14/MP0_IBNDR0/pmos_boundary
flabel space 20016 3024 20160 4032 0 FreeSans 320 90 0 0 I14/MP0_IBNDL0/pmos_boundary
flabel metal1 19986 2304 20046 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[0]/S0
flabel metal1 19842 2304 19902 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[0]/D0
flabel metal1 19698 2304 19758 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[0]/S1
flabel metal1 19786 2700 19960 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[0]/G0
rlabel pwell 20026 2670 20056 2692 1 I14/MN0_IM0[0]/BODY
flabel metal1 19698 2304 19758 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[1]/S0
flabel metal1 19554 2304 19614 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[1]/D0
flabel metal1 19410 2304 19470 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[1]/S1
flabel metal1 19498 2700 19672 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[1]/G0
rlabel pwell 19738 2670 19768 2692 1 I14/MN0_IM0[1]/BODY
flabel metal1 19410 2304 19470 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[2]/S0
flabel metal1 19266 2304 19326 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[2]/D0
flabel metal1 19122 2304 19182 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[2]/S1
flabel metal1 19210 2700 19384 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[2]/G0
rlabel pwell 19450 2670 19480 2692 1 I14/MN0_IM0[2]/BODY
flabel metal1 19122 2304 19182 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[3]/S0
flabel metal1 18978 2304 19038 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[3]/D0
flabel metal1 18834 2304 18894 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[3]/S1
flabel metal1 18922 2700 19096 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[3]/G0
rlabel pwell 19162 2670 19192 2692 1 I14/MN0_IM0[3]/BODY
flabel metal1 18834 2304 18894 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[4]/S0
flabel metal1 18690 2304 18750 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[4]/D0
flabel metal1 18546 2304 18606 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[4]/S1
flabel metal1 18634 2700 18808 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[4]/G0
rlabel pwell 18874 2670 18904 2692 1 I14/MN0_IM0[4]/BODY
flabel metal1 18546 2304 18606 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[5]/S0
flabel metal1 18402 2304 18462 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[5]/D0
flabel metal1 18258 2304 18318 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[5]/S1
flabel metal1 18346 2700 18520 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[5]/G0
rlabel pwell 18586 2670 18616 2692 1 I14/MN0_IM0[5]/BODY
flabel metal1 18258 2304 18318 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[6]/S0
flabel metal1 18114 2304 18174 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[6]/D0
flabel metal1 17970 2304 18030 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[6]/S1
flabel metal1 18058 2700 18232 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[6]/G0
rlabel pwell 18298 2670 18328 2692 1 I14/MN0_IM0[6]/BODY
flabel metal1 17970 2304 18030 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[7]/S0
flabel metal1 17826 2304 17886 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[7]/D0
flabel metal1 17682 2304 17742 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[7]/S1
flabel metal1 17770 2700 17944 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[7]/G0
rlabel pwell 18010 2670 18040 2692 1 I14/MN0_IM0[7]/BODY
flabel metal1 17682 2304 17742 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[8]/S0
flabel metal1 17538 2304 17598 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[8]/D0
flabel metal1 17394 2304 17454 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[8]/S1
flabel metal1 17482 2700 17656 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[8]/G0
rlabel pwell 17722 2670 17752 2692 1 I14/MN0_IM0[8]/BODY
flabel metal1 17394 2304 17454 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[9]/S0
flabel metal1 17250 2304 17310 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[9]/D0
flabel metal1 17106 2304 17166 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[9]/S1
flabel metal1 17194 2700 17368 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[9]/G0
rlabel pwell 17434 2670 17464 2692 1 I14/MN0_IM0[9]/BODY
flabel metal1 17106 2304 17166 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[10]/S0
flabel metal1 16962 2304 17022 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[10]/D0
flabel metal1 16818 2304 16878 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[10]/S1
flabel metal1 16906 2700 17080 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[10]/G0
rlabel pwell 17146 2670 17176 2692 1 I14/MN0_IM0[10]/BODY
flabel metal1 16818 2304 16878 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[11]/S0
flabel metal1 16674 2304 16734 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[11]/D0
flabel metal1 16530 2304 16590 2630 0 FreeSans 240 0 0 0 I14/MN0_IM0[11]/S1
flabel metal1 16618 2700 16792 2772 0 FreeSans 240 0 0 0 I14/MN0_IM0[11]/G0
rlabel pwell 16858 2670 16888 2692 1 I14/MN0_IM0[11]/BODY
flabel space 16416 2016 16560 3024 0 FreeSans 320 90 0 0 I14/MN0_IBNDR0/nmos_boundary
flabel space 20016 2016 20160 3024 0 FreeSans 320 90 0 0 I14/MN0_IBNDL0/nmos_boundary
flabel space 20160 3024 20304 4032 0 FreeSans 320 90 0 0 SPACE0[0]/pspace/PMOS_SPACE
flabel space 20160 2016 20304 3024 0 FreeSans 320 90 0 0 SPACE0[0]/nspace/NMOS_SPACE
flabel space 20304 3024 20448 4032 0 FreeSans 320 90 0 0 SPACE0[1]/pspace/PMOS_SPACE
flabel space 20304 2016 20448 3024 0 FreeSans 320 90 0 0 SPACE0[1]/nspace/NMOS_SPACE
flabel space 20448 3024 20592 4032 0 FreeSans 320 90 0 0 SPACE0[2]/pspace/PMOS_SPACE
flabel space 20448 2016 20592 3024 0 FreeSans 320 90 0 0 SPACE0[2]/nspace/NMOS_SPACE
flabel space 20592 3024 20736 4032 0 FreeSans 320 90 0 0 SPACE0[3]/pspace/PMOS_SPACE
flabel space 20592 2016 20736 3024 0 FreeSans 320 90 0 0 SPACE0[3]/nspace/NMOS_SPACE
flabel space 20736 3024 20880 4032 0 FreeSans 320 90 0 0 SPACE0[4]/pspace/PMOS_SPACE
flabel space 20736 2016 20880 3024 0 FreeSans 320 90 0 0 SPACE0[4]/nspace/NMOS_SPACE
flabel space 20880 3024 21024 4032 0 FreeSans 320 90 0 0 SPACE0[5]/pspace/PMOS_SPACE
flabel space 20880 2016 21024 3024 0 FreeSans 320 90 0 0 SPACE0[5]/nspace/NMOS_SPACE
<< end >>
