magic
tech sky130A
timestamp 1655825368
<< nwell >>
rect 0 66 72 342
<< labels >>
flabel space 0 0 72 504 0 FreeSans 160 90 0 0 PMOS_SPACE
<< end >>
