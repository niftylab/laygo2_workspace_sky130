magic
tech sky130A
timestamp 1679560919
<< checkpaint >>
rect -640 1638 928 1668
rect -640 -134 930 1638
rect -640 -660 928 -134
<< metal1 >>
rect 57 844 87 1028
rect 201 844 231 1028
rect 57 -20 87 164
rect 201 -20 231 164
<< metal2 >>
rect -10 978 298 1038
rect 72 777 216 807
rect 72 201 216 231
rect -10 -30 298 30
use ntap_fast_boundary  MNT0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825115
transform 1 0 0 0 1 0
box 0 0 72 512
use ntap_fast_boundary  MNT0_IBNDR0
timestamp 1655825115
transform 1 0 216 0 1 0
box 0 0 72 512
use ntap_fast_center_nf2_v2  MNT0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656694979
transform 1 0 72 0 1 0
box -36 143 180 342
use via_M1_M2_0  MNT0_IVTAP10 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 144 0 1 216
box -16 -16 16 16
use via_M1_M2_1  MNT0_IVTIETAP10 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 72 0 1 0
box -16 -16 16 16
use ptap_fast_boundary  MPT0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825477
transform 1 0 0 0 -1 1008
box 0 0 84 512
use ptap_fast_boundary  MPT0_IBNDR0
timestamp 1655825477
transform 1 0 216 0 -1 1008
box 0 0 84 512
use ptap_fast_center_nf2_v2  MPT0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656699071
transform 1 0 72 0 -1 1008
box -36 66 180 342
use via_M1_M2_0  MPT0_IVTAP10
timestamp 1647525606
transform 1 0 144 0 -1 792
box -16 -16 16 16
use via_M1_M2_1  MPT0_IVTIETAP10
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 72 0 -1 1008
box -16 -16 16 16
<< end >>
