magic
tech sky130A
timestamp 1655825115
<< pwell >>
rect 0 186 72 342
<< labels >>
flabel space 0 0 72 512 0 FreeSans 160 90 0 0 ntap_boundary
<< end >>
