magic
tech sky130A
magscale 1 2
timestamp 1704392934
<< locali >>
rect -17 -17 17 17
<< end >>
