magic
tech sky130A
timestamp 1679561080
<< checkpaint >>
rect -650 -660 38666 1668
<< metal2 >>
rect -20 978 38036 1038
rect 417 489 663 519
rect 705 489 1599 519
rect 7761 489 8079 519
rect 8337 489 8583 519
rect 11937 489 12255 519
rect 12513 489 12759 519
rect 16113 489 16431 519
rect 16689 489 16935 519
rect 20289 489 20607 519
rect 20865 489 21111 519
rect 24465 489 24783 519
rect 25041 489 25287 519
rect 28641 489 28959 519
rect 29217 489 29463 519
rect 32817 489 33135 519
rect 33393 489 33639 519
rect 36993 489 37311 519
rect 37569 489 37815 519
rect -20 -30 38036 30
<< metal3 >>
rect 129 129 159 375
rect 345 360 375 648
rect 417 129 447 519
rect 633 345 663 519
rect 705 201 735 519
rect 921 129 951 375
rect 1209 360 1239 648
rect 1569 345 1599 519
rect 993 201 1023 303
rect 4665 201 4695 375
rect 5313 360 5343 648
rect 7761 201 7791 519
rect 8049 345 8079 519
rect 8265 273 8295 375
rect 8337 129 8367 519
rect 8409 129 8439 375
rect 8553 345 8583 519
rect 8625 216 8655 792
rect 8841 201 8871 375
rect 9489 360 9519 648
rect 11937 201 11967 519
rect 12225 345 12255 519
rect 12441 273 12471 375
rect 12513 129 12543 519
rect 12585 129 12615 375
rect 12729 345 12759 519
rect 12801 216 12831 792
rect 13017 201 13047 375
rect 13665 360 13695 648
rect 16113 201 16143 519
rect 16401 345 16431 519
rect 16617 273 16647 375
rect 16689 129 16719 519
rect 16761 129 16791 375
rect 16905 345 16935 519
rect 16977 216 17007 792
rect 17193 201 17223 375
rect 17841 360 17871 648
rect 20289 201 20319 519
rect 20577 345 20607 519
rect 20793 273 20823 375
rect 20865 129 20895 519
rect 20937 129 20967 375
rect 21081 345 21111 519
rect 21153 216 21183 792
rect 21369 201 21399 375
rect 22017 360 22047 648
rect 24465 201 24495 519
rect 24753 345 24783 519
rect 24969 273 24999 375
rect 25041 129 25071 519
rect 25113 129 25143 375
rect 25257 345 25287 519
rect 25329 216 25359 792
rect 25545 201 25575 375
rect 26193 360 26223 648
rect 28641 201 28671 519
rect 28929 345 28959 519
rect 29145 273 29175 375
rect 29217 129 29247 519
rect 29289 129 29319 375
rect 29433 345 29463 519
rect 29505 216 29535 792
rect 29721 201 29751 375
rect 30369 360 30399 648
rect 32817 201 32847 519
rect 33105 345 33135 519
rect 33321 273 33351 375
rect 33393 129 33423 519
rect 33465 129 33495 375
rect 33609 345 33639 519
rect 33681 216 33711 792
rect 33897 201 33927 375
rect 34545 360 34575 648
rect 36993 201 37023 519
rect 37281 345 37311 519
rect 37497 273 37527 375
rect 37569 129 37599 519
rect 37641 129 37671 375
rect 37785 345 37815 519
rect 37857 216 37887 792
<< metal4 >>
rect 993 273 37527 303
rect 4449 201 33927 231
rect 129 129 37671 159
use logic_advanced_cgate_2x  cgate0 magic_layout/logic_advanced
timestamp 1679561063
transform 1 0 1152 0 1 0
box -20 -30 3476 1038
use logic_generated_dff_2x  dff_0 magic_layout/logic_generated
timestamp 1679561001
transform 1 0 4608 0 1 0
box -20 -30 3332 1038
use logic_generated_dff_2x  dff_1
timestamp 1679561001
transform 1 0 8784 0 1 0
box -20 -30 3332 1038
use logic_generated_dff_2x  dff_2
timestamp 1679561001
transform 1 0 12960 0 1 0
box -20 -30 3332 1038
use logic_generated_dff_2x  dff_3
timestamp 1679561001
transform 1 0 17136 0 1 0
box -20 -30 3332 1038
use logic_generated_dff_2x  dff_4
timestamp 1679561001
transform 1 0 21312 0 1 0
box -20 -30 3332 1038
use logic_generated_dff_2x  dff_5
timestamp 1679561001
transform 1 0 25488 0 1 0
box -20 -30 3332 1038
use logic_generated_dff_2x  dff_6
timestamp 1679561001
transform 1 0 29664 0 1 0
box -20 -30 3332 1038
use logic_generated_dff_2x  dff_7
timestamp 1679561001
transform 1 0 33840 0 1 0
box -20 -30 3332 1038
use logic_generated_inv_2x  inv0 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 8496 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv1
timestamp 1679560816
transform 1 0 12672 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv2
timestamp 1679560816
transform 1 0 16848 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv3
timestamp 1679560816
transform 1 0 21024 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv4
timestamp 1679560816
transform 1 0 25200 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv5
timestamp 1679560816
transform 1 0 29376 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv6
timestamp 1679560816
transform 1 0 33552 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv7
timestamp 1679560816
transform 1 0 37728 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv_and
timestamp 1679560816
transform 1 0 576 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv_sel
timestamp 1679560816
transform 1 0 864 0 1 0
box -20 -30 308 1038
use logic_generated_nand_2x  nand magic_layout/logic_generated
timestamp 1679560872
transform 1 0 0 0 1 0
box -20 -30 596 1038
use via_M3_M4_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 144 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_3
timestamp 1647526059
transform 1 0 936 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_5
timestamp 1647526059
transform 1 0 8424 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_7
timestamp 1647526059
transform 1 0 12600 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_9
timestamp 1647526059
transform 1 0 16776 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_11
timestamp 1647526059
transform 1 0 20952 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_13
timestamp 1647526059
transform 1 0 25128 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_15
timestamp 1647526059
transform 1 0 29304 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_17
timestamp 1647526059
transform 1 0 33480 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_19
timestamp 1647526059
transform 1 0 37656 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_22
timestamp 1647526059
transform 1 0 1008 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_24
timestamp 1647526059
transform 1 0 8280 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_26
timestamp 1647526059
transform 1 0 12456 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_28
timestamp 1647526059
transform 1 0 16632 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_30
timestamp 1647526059
transform 1 0 20808 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_32
timestamp 1647526059
transform 1 0 24984 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_34
timestamp 1647526059
transform 1 0 29160 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_36
timestamp 1647526059
transform 1 0 33336 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_38
timestamp 1647526059
transform 1 0 37512 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_41 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 432 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_43
timestamp 1647525786
transform 1 0 648 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_46
timestamp 1647525786
transform 1 0 720 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_48
timestamp 1647525786
transform 1 0 1584 0 1 504
box -19 -19 19 19
use via_M3_M4_0  NoName_50
timestamp 1647526059
transform 1 0 4464 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_52
timestamp 1647526059
transform 1 0 4680 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_54
timestamp 1647526059
transform 1 0 8856 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_56
timestamp 1647526059
transform 1 0 13032 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_58
timestamp 1647526059
transform 1 0 17208 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_60
timestamp 1647526059
transform 1 0 21384 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_62
timestamp 1647526059
transform 1 0 25560 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_64
timestamp 1647526059
transform 1 0 29736 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_66
timestamp 1647526059
transform 1 0 33912 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_69
timestamp 1647525786
transform 1 0 7776 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_71
timestamp 1647525786
transform 1 0 8064 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_74
timestamp 1647525786
transform 1 0 8352 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_76
timestamp 1647525786
transform 1 0 8568 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_79
timestamp 1647525786
transform 1 0 11952 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_81
timestamp 1647525786
transform 1 0 12240 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_84
timestamp 1647525786
transform 1 0 12528 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_86
timestamp 1647525786
transform 1 0 12744 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_89
timestamp 1647525786
transform 1 0 16128 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_91
timestamp 1647525786
transform 1 0 16416 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_94
timestamp 1647525786
transform 1 0 16704 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_96
timestamp 1647525786
transform 1 0 16920 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_99
timestamp 1647525786
transform 1 0 20304 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_101
timestamp 1647525786
transform 1 0 20592 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_104
timestamp 1647525786
transform 1 0 20880 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_106
timestamp 1647525786
transform 1 0 21096 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_109
timestamp 1647525786
transform 1 0 24480 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_111
timestamp 1647525786
transform 1 0 24768 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_114
timestamp 1647525786
transform 1 0 25056 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_116
timestamp 1647525786
transform 1 0 25272 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_119
timestamp 1647525786
transform 1 0 28656 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_121
timestamp 1647525786
transform 1 0 28944 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_124
timestamp 1647525786
transform 1 0 29232 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_126
timestamp 1647525786
transform 1 0 29448 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_129
timestamp 1647525786
transform 1 0 32832 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_131
timestamp 1647525786
transform 1 0 33120 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_134
timestamp 1647525786
transform 1 0 33408 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_136
timestamp 1647525786
transform 1 0 33624 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_139
timestamp 1647525786
transform 1 0 37008 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_141
timestamp 1647525786
transform 1 0 37296 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_144
timestamp 1647525786
transform 1 0 37584 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_146
timestamp 1647525786
transform 1 0 37800 0 1 504
box -19 -19 19 19
use logic_generated_tinv_2x  tinv0 magic_layout/logic_generated
timestamp 1679560906
transform 1 0 7920 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv1
timestamp 1679560906
transform 1 0 12096 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv2
timestamp 1679560906
transform 1 0 16272 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv3
timestamp 1679560906
transform 1 0 20448 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv4
timestamp 1679560906
transform 1 0 24624 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv5
timestamp 1679560906
transform 1 0 28800 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv6
timestamp 1679560906
transform 1 0 32976 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv7
timestamp 1679560906
transform 1 0 37152 0 1 0
box -20 -30 596 1038
<< labels >>
flabel metal3 1224 504 1224 504 0 FreeSans 240 90 0 0 CLK
port 1 nsew
flabel metal3 5328 504 5328 504 0 FreeSans 240 90 0 0 Di<0>
port 2 nsew
flabel metal3 9504 504 9504 504 0 FreeSans 240 90 0 0 Di<1>
port 3 nsew
flabel metal3 13680 504 13680 504 0 FreeSans 240 90 0 0 Di<2>
port 4 nsew
flabel metal3 17856 504 17856 504 0 FreeSans 240 90 0 0 Di<3>
port 5 nsew
flabel metal3 22032 504 22032 504 0 FreeSans 240 90 0 0 Di<4>
port 6 nsew
flabel metal3 26208 504 26208 504 0 FreeSans 240 90 0 0 Di<5>
port 7 nsew
flabel metal3 30384 504 30384 504 0 FreeSans 240 90 0 0 Di<6>
port 8 nsew
flabel metal3 34560 504 34560 504 0 FreeSans 240 90 0 0 Di<7>
port 9 nsew
flabel metal3 8640 504 8640 504 0 FreeSans 240 90 0 0 Do<0>
port 10 nsew
flabel metal3 12816 504 12816 504 0 FreeSans 240 90 0 0 Do<1>
port 11 nsew
flabel metal3 16992 504 16992 504 0 FreeSans 240 90 0 0 Do<2>
port 12 nsew
flabel metal3 21168 504 21168 504 0 FreeSans 240 90 0 0 Do<3>
port 13 nsew
flabel metal3 25344 504 25344 504 0 FreeSans 240 90 0 0 Do<4>
port 14 nsew
flabel metal3 29520 504 29520 504 0 FreeSans 240 90 0 0 Do<5>
port 15 nsew
flabel metal3 33696 504 33696 504 0 FreeSans 240 90 0 0 Do<6>
port 16 nsew
flabel metal3 37872 504 37872 504 0 FreeSans 240 90 0 0 Do<7>
port 17 nsew
flabel metal4 18900 144 18900 144 0 FreeSans 240 0 0 0 SEL
port 18 nsew
flabel metal2 19008 1008 19008 1008 0 FreeSans 480 0 0 0 VDD
port 19 nsew
flabel metal2 19008 0 19008 0 0 FreeSans 480 0 0 0 VSS
port 20 nsew
flabel metal3 360 504 360 504 0 FreeSans 240 90 0 0 WE
port 21 nsew
<< end >>
