magic
tech sky130A
timestamp 1656694979
<< pwell >>
rect -36 186 180 342
<< psubdiff >>
rect -15 286 159 307
rect -15 242 -10 286
rect 10 242 62 286
rect 82 242 134 286
rect 154 242 159 286
rect -15 221 159 242
<< psubdiffcont >>
rect -10 242 10 286
rect 62 242 82 286
rect 134 242 154 286
<< locali >>
rect -15 286 15 307
rect -15 242 -10 286
rect 10 242 15 286
rect -15 221 15 242
rect 57 286 87 307
rect 57 242 62 286
rect 82 242 87 286
rect 57 221 87 242
rect 129 286 159 307
rect 129 242 134 286
rect 154 242 159 286
rect 129 221 159 242
<< viali >>
rect -10 242 10 286
rect 62 242 82 286
rect 134 242 154 286
<< metal1 >>
rect -15 286 15 307
rect -15 242 -10 286
rect 10 242 15 286
rect -15 143 15 242
rect 57 286 87 307
rect 57 242 62 286
rect 82 242 87 286
rect 57 143 87 242
rect 129 286 159 307
rect 129 242 134 286
rect 154 242 159 286
rect 129 143 159 242
<< end >>
