magic
tech sky130A
timestamp 1679560883
<< checkpaint >>
rect -650 -660 1226 1668
<< metal1 >>
rect 57 844 87 1028
rect 201 844 231 1028
rect 57 -20 87 164
rect 201 -20 231 164
rect 345 -20 375 164
rect 489 -20 519 164
<< metal2 >>
rect -20 978 596 1038
rect 342 849 522 879
rect 54 777 542 807
rect 54 633 234 663
rect 342 633 522 663
rect 54 345 234 375
rect 342 345 522 375
rect 54 201 522 231
rect -20 -30 596 30
<< metal3 >>
rect 129 345 159 663
rect 345 345 375 663
rect 417 201 447 879
use nmos13_fast_boundary  MN0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 216 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654175211
transform 1 0 72 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN0_IVD0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 144 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN0_IVG0
timestamp 1647525606
transform 1 0 144 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN0_IVTIED0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 72 0 1 0
box -16 -16 16 16
use nmos13_fast_boundary  MN1_IBNDL0
timestamp 1655824928
transform 1 0 288 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN1_IBNDR0
timestamp 1655824928
transform 1 0 504 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN1_IM0
timestamp 1654175211
transform 1 0 360 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN1_IVD0
timestamp 1647525606
transform 1 0 432 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN1_IVG0
timestamp 1647525606
transform 1 0 432 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN1_IVTIED0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 360 0 1 0
box -16 -16 16 16
use pmos13_fast_boundary  MP0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 216 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654091791
transform 1 0 72 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP0_IVD0
timestamp 1647525606
transform 1 0 144 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP0_IVG0
timestamp 1647525606
transform 1 0 144 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP0_IVTIED0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 72 0 -1 1008
box -16 -16 16 16
use pmos13_fast_boundary  MP1_IBNDL0
timestamp 1655825313
transform 1 0 288 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP1_IBNDR0
timestamp 1655825313
transform 1 0 504 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP1_IM0
timestamp 1654091791
transform 1 0 360 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP1_IVD0
timestamp 1647525606
transform 1 0 432 0 -1 864
box -16 -16 16 16
use via_M1_M2_0  MP1_IVG0
timestamp 1647525606
transform 1 0 432 0 -1 648
box -16 -16 16 16
use via_M1_M2_0  MP1_IVS0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 360 0 -1 792
box -16 -16 16 16
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 360 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 360 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 144 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 144 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_10
timestamp 1647525786
transform 1 0 432 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_12
timestamp 1647525786
transform 1 0 432 0 1 864
box -19 -19 19 19
<< labels >>
flabel metal3 360 504 360 504 0 FreeSans 240 90 0 0 A
port 1 nsew
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 B
port 2 nsew
flabel metal3 432 540 432 540 0 FreeSans 240 90 0 0 OUT
port 3 nsew
flabel metal2 288 1008 288 1008 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel metal2 288 0 288 0 0 FreeSans 480 0 0 0 VSS
port 5 nsew
<< end >>
