magic
tech sky130A
timestamp 1679560937
<< checkpaint >>
rect -630 -630 702 1638
use nmos13_fast_space_1x  nspace ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825027
transform 1 0 0 0 1 0
box 0 0 72 504
use pmos13_fast_space_1x  pspace ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825383
transform 1 0 0 0 -1 1008
box 0 0 72 504
<< end >>
