magic
tech sky130A
timestamp 1679560990
<< checkpaint >>
rect -650 -660 2658 1668
<< metal1 >>
rect 57 844 87 1028
rect 201 844 231 1028
rect 1209 844 1239 1028
rect 1353 844 1383 1028
rect 1497 844 1527 1028
rect 1641 844 1671 1028
rect 57 -20 87 164
rect 201 -20 231 164
rect 1209 -20 1239 164
rect 1353 -20 1383 164
rect 1497 -20 1527 164
rect 1641 -20 1671 164
<< metal2 >>
rect -20 978 1748 1038
rect 322 849 1450 879
rect 54 777 522 807
rect 566 777 874 807
rect 918 777 1386 807
rect 1494 777 1674 807
rect 54 633 234 663
rect 342 633 586 663
rect 710 633 1098 663
rect 1206 633 1386 663
rect 1430 633 1674 663
rect 54 345 234 375
rect 342 345 730 375
rect 854 345 1098 375
rect 1206 345 1386 375
rect 1430 345 1674 375
rect 54 201 522 231
rect 918 201 1386 231
rect 1494 201 1674 231
rect 322 129 1118 159
rect -20 -30 1748 30
<< metal3 >>
rect 129 345 159 663
rect 561 633 591 879
rect 705 345 735 663
rect 849 345 879 807
rect 1065 129 1095 879
rect 1281 345 1311 663
rect 1425 345 1455 879
rect 1569 201 1599 807
use nmos13_fast_boundary  MN0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 216 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654175211
transform 1 0 72 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN0_IVD0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 144 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN0_IVG0
timestamp 1647525606
transform 1 0 144 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN0_IVTIED0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 72 0 1 0
box -16 -16 16 16
use nmos13_fast_boundary  MN1_IBNDL0
timestamp 1655824928
transform 1 0 288 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN1_IBNDR0
timestamp 1655824928
transform 1 0 504 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN1_IM0
timestamp 1654175211
transform 1 0 360 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN1_IVD0
timestamp 1647525606
transform 1 0 432 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN1_IVG0
timestamp 1647525606
transform 1 0 432 0 1 360
box -16 -16 16 16
use via_M1_M2_0  MN1_IVS0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 360 0 1 144
box -16 -16 16 16
use nmos13_fast_boundary  MN2_IBNDL0
timestamp 1655824928
transform 1 0 864 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN2_IBNDR0
timestamp 1655824928
transform 1 0 1080 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN2_IM0
timestamp 1654175211
transform 1 0 936 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN2_IVD0
timestamp 1647525606
transform 1 0 1008 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN2_IVG0
timestamp 1647525606
transform 1 0 1008 0 1 360
box -16 -16 16 16
use via_M1_M2_0  MN2_IVS0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 936 0 1 144
box -16 -16 16 16
use nmos13_fast_boundary  MN3_IBNDL0
timestamp 1655824928
transform 1 0 1152 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN3_IBNDR0
timestamp 1655824928
transform 1 0 1368 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN3_IM0
timestamp 1654175211
transform 1 0 1224 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN3_IVD0
timestamp 1647525606
transform 1 0 1296 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN3_IVG0
timestamp 1647525606
transform 1 0 1296 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN3_IVTIED0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 1224 0 1 0
box -16 -16 16 16
use nmos13_fast_boundary  MN4_IBNDL0
timestamp 1655824928
transform 1 0 1440 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN4_IBNDR0
timestamp 1655824928
transform 1 0 1656 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN4_IM0
timestamp 1654175211
transform 1 0 1512 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN4_IVD0
timestamp 1647525606
transform 1 0 1584 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN4_IVG0
timestamp 1647525606
transform 1 0 1584 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN4_IVTIED0
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 1512 0 1 0
box -16 -16 16 16
use pmos13_fast_boundary  MP0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 216 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654091791
transform 1 0 72 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP0_IVD0
timestamp 1647525606
transform 1 0 144 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP0_IVG0
timestamp 1647525606
transform 1 0 144 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP0_IVTIED0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 72 0 -1 1008
box -16 -16 16 16
use pmos13_fast_boundary  MP1_IBNDL0
timestamp 1655825313
transform 1 0 288 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP1_IBNDR0
timestamp 1655825313
transform 1 0 504 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP1_IM0
timestamp 1654091791
transform 1 0 360 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP1_IVD0
timestamp 1647525606
transform 1 0 432 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP1_IVG0
timestamp 1647525606
transform 1 0 432 0 -1 648
box -16 -16 16 16
use via_M1_M2_0  MP1_IVS0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 360 0 -1 864
box -16 -16 16 16
use pmos13_fast_boundary  MP2_IBNDL0
timestamp 1655825313
transform 1 0 864 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP2_IBNDR0
timestamp 1655825313
transform 1 0 1080 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP2_IM0
timestamp 1654091791
transform 1 0 936 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP2_IVD0
timestamp 1647525606
transform 1 0 1008 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP2_IVG0
timestamp 1647525606
transform 1 0 1008 0 -1 648
box -16 -16 16 16
use via_M1_M2_0  MP2_IVS0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 936 0 -1 864
box -16 -16 16 16
use pmos13_fast_boundary  MP3_IBNDL0
timestamp 1655825313
transform 1 0 1152 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP3_IBNDR0
timestamp 1655825313
transform 1 0 1368 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP3_IM0
timestamp 1654091791
transform 1 0 1224 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP3_IVD0
timestamp 1647525606
transform 1 0 1296 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP3_IVG0
timestamp 1647525606
transform 1 0 1296 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP3_IVTIED0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 1224 0 -1 1008
box -16 -16 16 16
use pmos13_fast_boundary  MP4_IBNDL0
timestamp 1655825313
transform 1 0 1440 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP4_IBNDR0
timestamp 1655825313
transform 1 0 1656 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP4_IM0
timestamp 1654091791
transform 1 0 1512 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP4_IVD0
timestamp 1647525606
transform 1 0 1584 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP4_IVG0
timestamp 1647525606
transform 1 0 1584 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP4_IVTIED0
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 1512 0 -1 1008
box -16 -16 16 16
use via_M2_M3_0  NoName_0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 144 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_2
timestamp 1647525786
transform 1 0 144 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 1296 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 1296 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_6
timestamp 1647525786
transform 1 0 1584 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_8
timestamp 1647525786
transform 1 0 1584 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_10
timestamp 1647525786
transform 1 0 720 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_12
timestamp 1647525786
transform 1 0 720 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_15
timestamp 1647525786
transform 1 0 864 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_17
timestamp 1647525786
transform 1 0 864 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_20
timestamp 1647525786
transform 1 0 576 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_21
timestamp 1647525786
transform 1 0 576 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_27
timestamp 1647525786
transform 1 0 1080 0 1 144
box -19 -19 19 19
use via_M2_M3_0  NoName_28
timestamp 1647525786
transform 1 0 1080 0 1 864
box -19 -19 19 19
use via_M2_M3_0  NoName_31
timestamp 1647525786
transform 1 0 1440 0 1 864
box -19 -19 19 19
use via_M2_M3_0  NoName_33
timestamp 1647525786
transform 1 0 1440 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_36
timestamp 1647525786
transform 1 0 1440 0 1 648
box -19 -19 19 19
use nmos13_fast_space_2x  nspace0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825056
transform 1 0 576 0 1 0
box 0 0 144 504
use nmos13_fast_space_2x  nspace1
timestamp 1655825056
transform 1 0 720 0 1 0
box 0 0 144 504
use pmos13_fast_space_2x  pspace0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825401
transform 1 0 576 0 -1 1008
box 0 0 144 504
use pmos13_fast_space_2x  pspace1
timestamp 1655825401
transform 1 0 720 0 -1 1008
box 0 0 144 504
use logic_generated_TAP  TAP0 magic_layout/logic_generated
timestamp 1679560919
transform 1 0 1728 0 1 0
box -10 -30 300 1038
<< labels >>
flabel metal3 720 504 720 504 0 FreeSans 240 90 0 0 EN0
port 1 nsew
flabel metal3 864 576 864 576 0 FreeSans 240 90 0 0 EN1
port 2 nsew
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 I0
port 3 nsew
flabel metal3 1296 504 1296 504 0 FreeSans 240 90 0 0 I1
port 4 nsew
flabel metal3 1584 504 1584 504 0 FreeSans 240 90 0 0 O
port 5 nsew
flabel metal2 864 1008 864 1008 0 FreeSans 480 0 0 0 VDD
port 6 nsew
flabel metal2 864 0 864 0 0 FreeSans 480 0 0 0 VSS
port 7 nsew
<< end >>
