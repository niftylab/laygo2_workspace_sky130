magic
tech sky130A
magscale 1 2
timestamp 1654175211
<< pwell >>
rect -92 372 380 684
<< nmoslvt >>
rect 56 408 86 648
rect 200 408 230 648
<< ndiff >>
rect -56 598 56 648
rect -56 558 -20 598
rect 20 558 56 598
rect -56 498 56 558
rect -56 458 -20 498
rect 20 458 56 498
rect -56 408 56 458
rect 86 598 200 648
rect 86 558 124 598
rect 164 558 200 598
rect 86 498 200 558
rect 86 458 124 498
rect 164 458 200 498
rect 86 408 200 458
rect 230 598 344 648
rect 230 558 268 598
rect 308 558 344 598
rect 230 498 344 558
rect 230 458 268 498
rect 308 458 344 498
rect 230 408 344 458
<< ndiffc >>
rect -20 558 20 598
rect -20 458 20 498
rect 124 558 164 598
rect 124 458 164 498
rect 268 558 308 598
rect 268 458 308 498
<< poly >>
rect 56 737 230 756
rect 56 703 76 737
rect 110 703 184 737
rect 218 703 230 737
rect 56 684 230 703
rect 56 648 86 684
rect 200 648 230 684
rect 56 372 86 408
rect 200 372 230 408
<< polycont >>
rect 76 703 110 737
rect 184 703 218 737
<< locali >>
rect 56 737 230 756
rect 56 703 76 737
rect 110 703 184 737
rect 218 703 230 737
rect 56 684 230 703
rect -30 598 30 614
rect -30 558 -20 598
rect 20 558 30 598
rect -30 498 30 558
rect -30 458 -20 498
rect 20 458 30 498
rect -30 442 30 458
rect 114 598 174 614
rect 114 558 124 598
rect 164 558 174 598
rect 114 498 174 558
rect 114 458 124 498
rect 164 458 174 498
rect 114 442 174 458
rect 258 598 318 614
rect 258 558 268 598
rect 308 558 318 598
rect 258 498 318 558
rect 258 458 268 498
rect 308 458 318 498
rect 258 442 318 458
<< viali >>
rect 76 703 110 737
rect 184 703 218 737
rect -20 558 20 598
rect -20 458 20 498
rect 124 558 164 598
rect 124 458 164 498
rect 268 558 308 598
rect 268 458 308 498
<< metal1 >>
rect 56 737 230 756
rect 56 703 76 737
rect 110 703 184 737
rect 218 703 230 737
rect 56 684 230 703
rect -30 598 30 614
rect -30 558 -20 598
rect 20 558 30 598
rect -30 498 30 558
rect -30 458 -20 498
rect 20 458 30 498
rect -30 286 30 458
rect 114 598 174 614
rect 114 558 124 598
rect 164 558 174 598
rect 114 498 174 558
rect 114 458 124 498
rect 164 458 174 498
rect 114 286 174 458
rect 258 598 318 614
rect 258 558 268 598
rect 308 558 318 598
rect 258 498 318 558
rect 258 458 268 498
rect 308 458 318 498
rect 258 286 318 458
<< labels >>
flabel metal1 -30 288 30 614 0 FreeSans 240 0 0 0 S0
port 3 nsew
flabel metal1 114 288 174 614 0 FreeSans 240 0 0 0 D0
port 1 nsew
flabel metal1 258 288 318 614 0 FreeSans 240 0 0 0 S1
port 4 nsew
flabel metal1 56 684 230 756 0 FreeSans 240 0 0 0 G0
port 2 nsew
rlabel pwell -40 654 -10 676 1 BODY
port 5 nsew
<< end >>
