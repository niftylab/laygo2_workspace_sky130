magic
tech sky130A
timestamp 1679560942
<< checkpaint >>
rect -650 -660 938 1668
<< metal2 >>
rect -20 978 308 1038
rect -20 -30 308 30
use nmos13_fast_space_1x  nspace ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 3 72 0 0 504
timestamp 1655825027
transform 1 0 0 0 1 0
box 0 0 72 504
use pmos13_fast_space_1x  pspace ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 3 72 0 0 -504
timestamp 1655825383
transform 1 0 0 0 -1 1008
box 0 0 72 504
<< labels >>
flabel metal2 144 1008 144 1008 0 FreeSans 480 0 0 0 VDD
port 1 nsew
flabel metal2 144 0 144 0 0 FreeSans 480 0 0 0 VSS
port 2 nsew
<< end >>
