** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/byte_dff.sch
.subckt byte_dff Di<7> Do<6> Di<6> Do<5> Di<5> Di<4> Do<3> Di<3> Do<2> Di<2> Do<1> Di<1> Do<0> Di<0>
+ WE SEL CLK VDD VSS Do<7> Do<4>
*.PININFO Di<7>:I Do<6>:O Di<6>:I Do<5>:O Di<5>:I Di<4>:I Do<3>:O Di<3>:I Do<2>:O Di<2>:I Do<1>:O
*+ Di<1>:I Do<0>:O Di<0>:I WE:I SEL:I CLK:I VDD:B VSS:B Do<7>:O Do<4>:O
X_nand1 SEL WE net2 VDD VSS nand NF=2
X_inv2 SEL VDD VSS SEL_bar inv NF=2
x1 VDD net3 ck_o CLK VSS clk_gate NF=2
xDFF1 VDD VSS Di<7> net18 ck_o DFF NF=2
X_inv1 net2 VDD VSS net3 inv NF=2
X_tinv0 net4 SEL SEL_bar VDD VSS Do<0> tinv NF=2
xDFF2 VDD VSS Di<6> net15 ck_o DFF NF=2
xDFF3 VDD VSS Di<5> net13 ck_o DFF NF=2
xDFF4 VDD VSS Di<4> net11 ck_o DFF NF=2
xDFF5 VDD VSS Di<3> net9 ck_o DFF NF=2
xDFF6 VDD VSS Di<2> net7 ck_o DFF NF=2
xDFF7 VDD VSS Di<1> net5 ck_o DFF NF=2
xDFF8 VDD VSS Di<0> net1 ck_o DFF NF=2
X_inv3 net1 VDD VSS net4 inv NF=2
X_tinv1 net6 SEL SEL_bar VDD VSS Do<1> tinv NF=2
X_inv4 net5 VDD VSS net6 inv NF=2
X_tinv2 net8 SEL SEL_bar VDD VSS Do<2> tinv NF=2
X_inv5 net7 VDD VSS net8 inv NF=2
X_tinv3 net10 SEL SEL_bar VDD VSS Do<3> tinv NF=2
X_inv6 net9 VDD VSS net10 inv NF=2
X_tinv4 net12 SEL SEL_bar VDD VSS Do<4> tinv NF=2
X_inv7 net11 VDD VSS net12 inv NF=2
X_tinv8 net14 SEL SEL_bar VDD VSS Do<5> tinv NF=2
X_inv9 net13 VDD VSS net14 inv NF=2
X_tinv10 net16 SEL SEL_bar VDD VSS Do<6> tinv NF=2
X_inv11 net15 VDD VSS net16 inv NF=2
X_tinv12 net17 SEL SEL_bar VDD VSS Do<7> tinv NF=2
X_inv13 net18 VDD VSS net17 inv NF=2
.ends

* expanding   symbol:  ./nand.sym # of pins=5
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nand.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nand.sch
.subckt nand B A Y VDD VSS  NF=2
*.PININFO Y:O A:I VDD:B VSS:B B:I
XM1 Y A net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM2 net1 B VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM3 Y B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
XM4 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
.ends


* expanding   symbol:  ./inv.sym # of pins=4
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/inv.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/inv.sch
.subckt inv X VDD VSS Y  NF=2
*.PININFO VSS:B X:I Y:O VDD:B
XM1 Y X VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM2 Y X VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
.ends


* expanding   symbol:  ./clk_gate.sym # of pins=5
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/clk_gate.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/clk_gate.sch
.subckt clk_gate VDD EN CK_O CK_I VSS  NF=2
*.PININFO CK_I:I VDD:B VSS:B EN:I CK_O:O
X_inv1 CK_I VDD VSS net1 inv NF=2
X_latch1 EN net1 CK_I VSS VDD net2 latch NF=2
X_nand1 CK_I net2 net3 VDD VSS nand NF=2
X_inv2 net3 VDD VSS CK_O inv NF=2
.ends


* expanding   symbol:  ./DFF.sym # of pins=5
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/DFF.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/DFF.sch
.subckt DFF VDD VSS I O CLK  NF=2
*.PININFO VDD:B VSS:B I:I CLK:I O:O
X_latch1 I clk_bar clk_buf VSS VDD net1 latch NF=2
X_latch2 net1 clk_buf clk_bar VSS VDD O latch NF=2
X_inv1 CLK VDD VSS clk_bar inv NF=2
X_inv2 clk_bar VDD VSS clk_buf inv NF=2
.ends


* expanding   symbol:  ./tinv.sym # of pins=6
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/tinv.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/tinv.sch
.subckt tinv X EN ENB VDD VSS Y  NF=2
*.PININFO X:I ENB:I EN:I Y:O VDD:B VSS:B
XM1 net2 X VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
XM2 Y ENB net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
XM3 Y EN net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM4 net1 X VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
.ends


* expanding   symbol:  latch.sym # of pins=6
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/latch.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/latch.sch
.subckt latch IN CLK CLKB VSS VDD OUT  NF=2
*.PININFO CLKB:I IN:I CLK:I VDD:B VSS:B OUT:O
X_tinv1 IN CLK CLKB VDD VSS net1 tinv NF=NF
X_inv1 net1 VDD VSS OUT inv NF=NF
X_tinv_small1 OUT CLKB CLK VDD VSS net1 tinv_small
.ends


* expanding   symbol:  tinv_small.sym # of pins=6
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/tinv_small.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/tinv_small.sch
.subckt tinv_small X EN ENB VDD VSS Y
*.PININFO X:I ENB:I EN:I Y:O VDD:B VSS:B
XM1 net2 X VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=1
XM2 Y ENB net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=1
XM3 Y EN net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=1
XM4 net1 X VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=1
.ends

.end
