magic
tech sky130A
timestamp 1704386328
<< locali >>
rect -13 10 13 13
rect -13 -13 13 -10
<< viali >>
rect -13 -10 13 10
<< metal1 >>
rect -13 10 13 13
rect -13 -13 13 -10
<< end >>
