magic
tech sky130A
timestamp 1679561084
<< checkpaint >>
rect -650 -660 156170 1668
<< metal2 >>
rect -20 978 155540 1038
rect -20 -30 155540 30
<< metal3 >>
rect 345 360 375 648
rect 5313 360 5343 648
rect 8625 216 8655 792
rect 9489 360 9519 648
rect 12801 216 12831 792
rect 13665 360 13695 648
rect 16977 216 17007 792
rect 17841 360 17871 648
rect 21153 216 21183 792
rect 22017 360 22047 648
rect 25329 216 25359 792
rect 26193 360 26223 648
rect 29505 216 29535 792
rect 30369 360 30399 648
rect 33681 216 33711 792
rect 34545 360 34575 648
rect 37857 216 37887 792
rect 129 57 159 159
rect 38073 57 38103 375
rect 38433 57 38463 231
rect 39009 201 39039 375
rect 39513 360 39543 648
rect 44481 360 44511 648
rect 47793 216 47823 792
rect 48657 360 48687 648
rect 51969 216 51999 792
rect 52833 360 52863 648
rect 56145 216 56175 792
rect 57009 360 57039 648
rect 60321 216 60351 792
rect 61185 360 61215 648
rect 64497 216 64527 792
rect 65361 360 65391 648
rect 68673 216 68703 792
rect 69537 360 69567 648
rect 72849 216 72879 792
rect 73713 360 73743 648
rect 77025 216 77055 792
rect 39297 57 39327 159
rect 77241 57 77271 375
rect 77601 57 77631 231
rect 78177 201 78207 375
rect 78681 360 78711 648
rect 83649 360 83679 648
rect 86961 216 86991 792
rect 87825 360 87855 648
rect 91137 216 91167 792
rect 92001 360 92031 648
rect 95313 216 95343 792
rect 96177 360 96207 648
rect 99489 216 99519 792
rect 100353 360 100383 648
rect 103665 216 103695 792
rect 104529 360 104559 648
rect 107841 216 107871 792
rect 108705 360 108735 648
rect 112017 216 112047 792
rect 112881 360 112911 648
rect 116193 216 116223 792
rect 78465 57 78495 159
rect 116409 57 116439 375
rect 116769 57 116799 231
rect 117345 201 117375 375
rect 117849 360 117879 648
rect 122817 360 122847 648
rect 126129 216 126159 792
rect 126993 360 127023 648
rect 130305 216 130335 792
rect 131169 360 131199 648
rect 134481 216 134511 792
rect 135345 360 135375 648
rect 138657 216 138687 792
rect 139521 360 139551 648
rect 142833 216 142863 792
rect 143697 360 143727 648
rect 147009 216 147039 792
rect 147873 360 147903 648
rect 151185 216 151215 792
rect 152049 360 152079 648
rect 155361 216 155391 792
rect 117633 57 117663 159
<< metal4 >>
rect 1209 345 38679 375
rect 39009 345 77847 375
rect 78177 345 117015 375
rect 117345 345 118743 375
rect 129 57 38103 87
rect 38433 57 77271 87
rect 77601 57 116439 87
rect 116769 57 117663 87
use logic_generated_buffer_2x  buf_ck0 magic_layout/logic_generated
timestamp 1679560840
transform 1 0 38592 0 1 0
box -20 -30 596 1038
use logic_generated_buffer_2x  buf_ck1
timestamp 1679560840
transform 1 0 77760 0 1 0
box -20 -30 596 1038
use logic_generated_buffer_2x  buf_ck2
timestamp 1679560840
transform 1 0 116928 0 1 0
box -20 -30 596 1038
use logic_generated_buffer_2x  buf_sel0
timestamp 1679560840
transform 1 0 38016 0 1 0
box -20 -30 596 1038
use logic_generated_buffer_2x  buf_sel1
timestamp 1679560840
transform 1 0 77184 0 1 0
box -20 -30 596 1038
use logic_generated_buffer_2x  buf_sel2
timestamp 1679560840
transform 1 0 116352 0 1 0
box -20 -30 596 1038
use logic_advanced_byte_dff_2x  byte_dff0 magic_layout/logic_advanced
timestamp 1679561080
transform 1 0 0 0 1 0
box -20 -30 38036 1038
use logic_advanced_byte_dff_2x  byte_dff1
timestamp 1679561080
transform 1 0 39168 0 1 0
box -20 -30 38036 1038
use logic_advanced_byte_dff_2x  byte_dff2
timestamp 1679561080
transform 1 0 78336 0 1 0
box -20 -30 38036 1038
use logic_advanced_byte_dff_2x  byte_dff3
timestamp 1679561080
transform 1 0 117504 0 1 0
box -20 -30 38036 1038
use via_M3_M4_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 144 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_3
timestamp 1647526059
transform 1 0 38088 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_6
timestamp 1647526059
transform 1 0 38448 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_8
timestamp 1647526059
transform 1 0 39312 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_13
timestamp 1647526059
transform 1 0 77256 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_16
timestamp 1647526059
transform 1 0 77616 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_18
timestamp 1647526059
transform 1 0 78480 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_23
timestamp 1647526059
transform 1 0 116424 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_26
timestamp 1647526059
transform 1 0 116784 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_28
timestamp 1647526059
transform 1 0 117648 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_30
timestamp 1647526059
transform 1 0 1224 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_31
timestamp 1647526059
transform 1 0 38664 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_34
timestamp 1647526059
transform 1 0 39024 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_35
timestamp 1647526059
transform 1 0 40392 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_38
timestamp 1647526059
transform 1 0 77832 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_41
timestamp 1647526059
transform 1 0 78192 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_42
timestamp 1647526059
transform 1 0 79560 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_45
timestamp 1647526059
transform 1 0 117000 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_48
timestamp 1647526059
transform 1 0 117360 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_49
timestamp 1647526059
transform 1 0 118728 0 1 360
box -19 -19 19 19
<< labels >>
flabel metal4 19944 360 19944 360 0 FreeSans 240 0 0 0 CLK
port 1 nsew
flabel metal3 152064 504 152064 504 0 FreeSans 240 90 0 0 Di<0>
port 2 nsew
flabel metal3 147888 504 147888 504 0 FreeSans 240 90 0 0 Di<1>
port 3 nsew
flabel metal3 143712 504 143712 504 0 FreeSans 240 90 0 0 Di<2>
port 4 nsew
flabel metal3 139536 504 139536 504 0 FreeSans 240 90 0 0 Di<3>
port 5 nsew
flabel metal3 135360 504 135360 504 0 FreeSans 240 90 0 0 Di<4>
port 6 nsew
flabel metal3 131184 504 131184 504 0 FreeSans 240 90 0 0 Di<5>
port 7 nsew
flabel metal3 127008 504 127008 504 0 FreeSans 240 90 0 0 Di<6>
port 8 nsew
flabel metal3 122832 504 122832 504 0 FreeSans 240 90 0 0 Di<7>
port 9 nsew
flabel metal3 112896 504 112896 504 0 FreeSans 240 90 0 0 Di<8>
port 10 nsew
flabel metal3 108720 504 108720 504 0 FreeSans 240 90 0 0 Di<9>
port 11 nsew
flabel metal3 104544 504 104544 504 0 FreeSans 240 90 0 0 Di<10>
port 12 nsew
flabel metal3 100368 504 100368 504 0 FreeSans 240 90 0 0 Di<11>
port 13 nsew
flabel metal3 96192 504 96192 504 0 FreeSans 240 90 0 0 Di<12>
port 14 nsew
flabel metal3 92016 504 92016 504 0 FreeSans 240 90 0 0 Di<13>
port 15 nsew
flabel metal3 87840 504 87840 504 0 FreeSans 240 90 0 0 Di<14>
port 16 nsew
flabel metal3 83664 504 83664 504 0 FreeSans 240 90 0 0 Di<15>
port 17 nsew
flabel metal3 73728 504 73728 504 0 FreeSans 240 90 0 0 Di<16>
port 18 nsew
flabel metal3 69552 504 69552 504 0 FreeSans 240 90 0 0 Di<17>
port 19 nsew
flabel metal3 65376 504 65376 504 0 FreeSans 240 90 0 0 Di<18>
port 20 nsew
flabel metal3 61200 504 61200 504 0 FreeSans 240 90 0 0 Di<19>
port 21 nsew
flabel metal3 57024 504 57024 504 0 FreeSans 240 90 0 0 Di<20>
port 22 nsew
flabel metal3 52848 504 52848 504 0 FreeSans 240 90 0 0 Di<21>
port 23 nsew
flabel metal3 48672 504 48672 504 0 FreeSans 240 90 0 0 Di<22>
port 24 nsew
flabel metal3 44496 504 44496 504 0 FreeSans 240 90 0 0 Di<23>
port 25 nsew
flabel metal3 34560 504 34560 504 0 FreeSans 240 90 0 0 Di<24>
port 26 nsew
flabel metal3 30384 504 30384 504 0 FreeSans 240 90 0 0 Di<25>
port 27 nsew
flabel metal3 26208 504 26208 504 0 FreeSans 240 90 0 0 Di<26>
port 28 nsew
flabel metal3 22032 504 22032 504 0 FreeSans 240 90 0 0 Di<27>
port 29 nsew
flabel metal3 17856 504 17856 504 0 FreeSans 240 90 0 0 Di<28>
port 30 nsew
flabel metal3 13680 504 13680 504 0 FreeSans 240 90 0 0 Di<29>
port 31 nsew
flabel metal3 9504 504 9504 504 0 FreeSans 240 90 0 0 Di<30>
port 32 nsew
flabel metal3 5328 504 5328 504 0 FreeSans 240 90 0 0 Di<31>
port 33 nsew
flabel metal3 155376 504 155376 504 0 FreeSans 240 90 0 0 Do<0>
port 34 nsew
flabel metal3 151200 504 151200 504 0 FreeSans 240 90 0 0 Do<1>
port 35 nsew
flabel metal3 147024 504 147024 504 0 FreeSans 240 90 0 0 Do<2>
port 36 nsew
flabel metal3 142848 504 142848 504 0 FreeSans 240 90 0 0 Do<3>
port 37 nsew
flabel metal3 138672 504 138672 504 0 FreeSans 240 90 0 0 Do<4>
port 38 nsew
flabel metal3 134496 504 134496 504 0 FreeSans 240 90 0 0 Do<5>
port 39 nsew
flabel metal3 130320 504 130320 504 0 FreeSans 240 90 0 0 Do<6>
port 40 nsew
flabel metal3 126144 504 126144 504 0 FreeSans 240 90 0 0 Do<7>
port 41 nsew
flabel metal3 116208 504 116208 504 0 FreeSans 240 90 0 0 Do<8>
port 42 nsew
flabel metal3 112032 504 112032 504 0 FreeSans 240 90 0 0 Do<9>
port 43 nsew
flabel metal3 107856 504 107856 504 0 FreeSans 240 90 0 0 Do<10>
port 44 nsew
flabel metal3 103680 504 103680 504 0 FreeSans 240 90 0 0 Do<11>
port 45 nsew
flabel metal3 99504 504 99504 504 0 FreeSans 240 90 0 0 Do<12>
port 46 nsew
flabel metal3 95328 504 95328 504 0 FreeSans 240 90 0 0 Do<13>
port 47 nsew
flabel metal3 91152 504 91152 504 0 FreeSans 240 90 0 0 Do<14>
port 48 nsew
flabel metal3 86976 504 86976 504 0 FreeSans 240 90 0 0 Do<15>
port 49 nsew
flabel metal3 77040 504 77040 504 0 FreeSans 240 90 0 0 Do<16>
port 50 nsew
flabel metal3 72864 504 72864 504 0 FreeSans 240 90 0 0 Do<17>
port 51 nsew
flabel metal3 68688 504 68688 504 0 FreeSans 240 90 0 0 Do<18>
port 52 nsew
flabel metal3 64512 504 64512 504 0 FreeSans 240 90 0 0 Do<19>
port 53 nsew
flabel metal3 60336 504 60336 504 0 FreeSans 240 90 0 0 Do<20>
port 54 nsew
flabel metal3 56160 504 56160 504 0 FreeSans 240 90 0 0 Do<21>
port 55 nsew
flabel metal3 51984 504 51984 504 0 FreeSans 240 90 0 0 Do<22>
port 56 nsew
flabel metal3 47808 504 47808 504 0 FreeSans 240 90 0 0 Do<23>
port 57 nsew
flabel metal3 37872 504 37872 504 0 FreeSans 240 90 0 0 Do<24>
port 58 nsew
flabel metal3 33696 504 33696 504 0 FreeSans 240 90 0 0 Do<25>
port 59 nsew
flabel metal3 29520 504 29520 504 0 FreeSans 240 90 0 0 Do<26>
port 60 nsew
flabel metal3 25344 504 25344 504 0 FreeSans 240 90 0 0 Do<27>
port 61 nsew
flabel metal3 21168 504 21168 504 0 FreeSans 240 90 0 0 Do<28>
port 62 nsew
flabel metal3 16992 504 16992 504 0 FreeSans 240 90 0 0 Do<29>
port 63 nsew
flabel metal3 12816 504 12816 504 0 FreeSans 240 90 0 0 Do<30>
port 64 nsew
flabel metal3 8640 504 8640 504 0 FreeSans 240 90 0 0 Do<31>
port 65 nsew
flabel metal4 19116 72 19116 72 0 FreeSans 240 0 0 0 SEL
port 66 nsew
flabel metal2 77760 1008 77760 1008 0 FreeSans 480 0 0 0 VDD
port 67 nsew
flabel metal2 77760 0 77760 0 0 FreeSans 480 0 0 0 VSS
port 68 nsew
flabel metal3 117864 504 117864 504 0 FreeSans 240 90 0 0 WE<0>
port 69 nsew
flabel metal3 78696 504 78696 504 0 FreeSans 240 90 0 0 WE<1>
port 70 nsew
flabel metal3 39528 504 39528 504 0 FreeSans 240 90 0 0 WE<2>
port 71 nsew
flabel metal3 360 504 360 504 0 FreeSans 240 90 0 0 WE<3>
port 72 nsew
<< end >>
