magic
tech sky130A
timestamp 1656699071
<< nwell >>
rect -36 66 180 342
<< nsubdiff >>
rect -15 240 159 252
rect -15 164 -10 240
rect 10 164 62 240
rect 82 164 134 240
rect 154 164 159 240
rect -15 152 159 164
<< nsubdiffcont >>
rect -10 164 10 240
rect 62 164 82 240
rect 134 164 154 240
<< locali >>
rect -15 240 15 252
rect -15 164 -10 240
rect 10 164 15 240
rect -15 152 15 164
rect 57 240 87 252
rect 57 164 62 240
rect 82 164 87 240
rect 57 152 87 164
rect 129 240 159 252
rect 129 164 134 240
rect 154 164 159 240
rect 129 152 159 164
<< viali >>
rect -10 164 10 240
rect 62 164 82 240
rect 134 164 154 240
<< metal1 >>
rect -15 240 15 252
rect -15 164 -10 240
rect 10 164 15 240
rect -15 94 15 164
rect 57 240 87 252
rect 57 164 62 240
rect 82 164 87 240
rect 57 94 87 164
rect 129 240 159 252
rect 129 164 134 240
rect 154 164 159 240
rect 129 94 159 164
<< end >>
