magic
tech sky130A
magscale 1 2
timestamp 1706255560
<< checkpaint >>
rect -1336 2174 11414 2986
rect -1336 -514 11456 2174
rect -1277 -1326 11456 -514
rect 8676 -2156 11456 -1326
<< error_s >>
rect 164 813 204 847
rect 532 813 572 847
rect 900 813 940 847
rect 8260 813 8300 847
rect 8628 813 8668 847
rect 8812 813 8852 847
rect 9180 813 9220 847
rect 9364 813 9404 847
rect 9548 813 9588 847
rect 9732 813 9772 847
<< locali >>
rect 627 1228 937 1262
rect 167 398 1305 432
rect 6791 398 7101 432
rect 7527 398 7837 432
<< metal1 >>
rect 152 1079 216 1411
rect 244 1053 308 1188
rect 612 1136 676 1271
rect 888 1053 952 1271
rect 980 1053 1044 1188
rect 1348 1162 1412 1328
rect 1532 1162 1596 1328
rect 1900 1053 1964 1188
rect 5672 1053 5736 1188
rect 6040 1053 6104 1354
rect 6408 1162 6472 1328
rect 7144 1162 7208 1328
rect 7328 1136 7392 1354
rect 8248 970 8312 1437
rect 8616 1079 8680 1411
rect 60 306 124 607
rect 152 223 216 441
rect 520 332 584 498
rect 1256 306 1320 441
rect 1440 223 1504 607
rect 1992 332 2056 498
rect 2360 223 2424 607
rect 3464 306 3528 607
rect 6408 223 6472 607
rect 6684 306 6748 607
rect 6776 223 6840 441
rect 7052 306 7116 441
rect 7144 223 7208 607
rect 7420 306 7484 607
rect 7512 223 7576 441
rect 7788 306 7852 441
rect 7880 249 7944 581
rect 8248 223 8312 524
rect 8340 306 8404 607
rect 8524 306 8588 524
rect 8800 223 8864 607
rect 9076 306 9140 607
<< metal2 >>
rect 5954 1302 7386 1354
rect 1354 1136 2234 1188
rect 2550 1136 2786 1188
rect 5678 1136 7938 1188
rect 9542 1136 10054 1188
rect 250 1053 578 1105
rect 986 1053 1314 1105
rect 1630 1053 1958 1105
rect 8070 970 8306 1022
rect 66 555 1498 607
rect 2366 555 3522 607
rect 6414 555 6742 607
rect 7150 555 7478 607
rect 8070 555 8398 607
rect 8806 555 9134 607
rect 9542 555 9778 607
rect 2182 472 2694 524
rect 8254 472 8582 524
rect 2550 389 6466 441
<< metal3 >>
rect 2164 469 2252 1191
rect 2532 386 2620 1191
rect 8052 552 8140 1025
rect 9524 552 9612 1191
use logic_ver2_space_1x  FILL /WORK/hjpark/laygo2_workspace_sky130/magic_layout/logic_ver2
array 0 1 92 0 0 -830
timestamp 1706176348
transform 1 0 9936 0 -1 830
box 0 -84 168 1726
use logic_ver2_inv_2x  I0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/logic_ver2
timestamp 1706249504
transform 1 0 0 0 -1 830
box -17 -84 444 896
use logic_ver2_mux2to1_2x  I1 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/logic_ver2
timestamp 1706249538
transform 1 0 368 0 -1 830
box -17 -84 2284 896
use logic_ver2_dff_2x  I2 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/logic_ver2
timestamp 1706249534
transform 1 0 2576 0 -1 830
box -17 -84 4124 896
use logic_ver2_inv_2x  I3
timestamp 1706249504
transform 1 0 5888 0 1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I4
timestamp 1706249504
transform 1 0 6624 0 -1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I5
timestamp 1706249504
transform 1 0 6992 0 -1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I6
timestamp 1706249504
transform 1 0 7360 0 -1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I7
timestamp 1706249504
transform 1 0 7728 0 -1 830
box -17 -84 444 896
use logic_ver2_inv_16x  I14 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/logic_ver2
timestamp 1706174759
transform -1 0 10120 0 1 830
box -34 -84 1732 896
use logic_ver2_inv_2x  I15
timestamp 1706249504
transform -1 0 368 0 1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I16
timestamp 1706249504
transform -1 0 736 0 1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I17
timestamp 1706249504
transform -1 0 1104 0 1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I18
timestamp 1706249504
transform -1 0 1472 0 1 830
box -17 -84 444 896
use logic_ver2_inv_2x  I19
timestamp 1706249504
transform 1 0 1472 0 1 830
box -17 -84 444 896
use logic_ver2_dff_2x  I20
timestamp 1706249534
transform 1 0 1840 0 1 830
box -17 -84 4124 896
use logic_ver2_mux2to1_2x  I21
timestamp 1706249538
transform 1 0 6256 0 1 830
box -17 -84 2284 896
use logic_ver2_inv_2x  I22
timestamp 1706249504
transform -1 0 8464 0 -1 830
box -17 -84 444 896
use logic_ver2_inv_4x  I23 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/logic_ver2
timestamp 1706249504
transform 1 0 8464 0 -1 830
box -17 -84 628 896
use logic_ver2_inv_8x  I24 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/logic_ver2
timestamp 1706176164
transform 1 0 9016 0 -1 830
box -34 -84 996 896
use via_M3_M4_0  NoName_1 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704387757
transform 1 0 92 0 1 581
box -32 -26 32 26
use via_M3_M4_0  NoName_3
timestamp 1704387757
transform 1 0 1472 0 1 581
box -32 -26 32 26
use via_M2_M3_0  NoName_6 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704386899
transform 1 0 184 0 1 415
box -32 -17 32 17
use via_M2_M3_0  NoName_8
timestamp 1704386899
transform 1 0 1288 0 1 415
box -32 -17 32 17
use via_M3_M4_0  NoName_11
timestamp 1704387757
transform 1 0 2392 0 1 581
box -32 -26 32 26
use via_M3_M4_0  NoName_13
timestamp 1704387757
transform 1 0 3496 0 1 581
box -32 -26 32 26
use via_M4_M5_0  NoName_16 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706182685
transform 1 0 2208 0 1 1162
box -37 -34 37 34
use via_M4_M5_0  NoName_18
timestamp 1706182685
transform 1 0 2208 0 1 498
box -37 -34 37 34
use via_M3_M4_0  NoName_20
timestamp 1704387757
transform 1 0 1380 0 1 1162
box -32 -26 32 26
use via_M3_M4_0  NoName_21
timestamp 1704387757
transform 1 0 2668 0 1 498
box -32 -26 32 26
use via_M3_M4_0  NoName_23
timestamp 1704387757
transform 1 0 6440 0 1 581
box -32 -26 32 26
use via_M3_M4_0  NoName_25
timestamp 1704387757
transform 1 0 6716 0 1 581
box -32 -26 32 26
use via_M2_M3_0  NoName_28
timestamp 1704386899
transform 1 0 6808 0 1 415
box -32 -17 32 17
use via_M2_M3_0  NoName_30
timestamp 1704386899
transform 1 0 7084 0 1 415
box -32 -17 32 17
use via_M3_M4_0  NoName_33
timestamp 1704387757
transform 1 0 7176 0 1 581
box -32 -26 32 26
use via_M3_M4_0  NoName_35
timestamp 1704387757
transform 1 0 7452 0 1 581
box -32 -26 32 26
use via_M2_M3_0  NoName_38
timestamp 1704386899
transform 1 0 7544 0 1 415
box -32 -17 32 17
use via_M2_M3_0  NoName_40
timestamp 1704386899
transform 1 0 7820 0 1 415
box -32 -17 32 17
use via_M3_M4_0  NoName_42
timestamp 1704387757
transform 1 0 1288 0 1 1079
box -32 -26 32 26
use via_M3_M4_0  NoName_44
timestamp 1704387757
transform 1 0 1012 0 1 1079
box -32 -26 32 26
use via_M2_M3_0  NoName_47
timestamp 1704386899
transform 1 0 920 0 1 1245
box -32 -17 32 17
use via_M2_M3_0  NoName_49
timestamp 1704386899
transform 1 0 644 0 1 1245
box -32 -17 32 17
use via_M3_M4_0  NoName_51
timestamp 1704387757
transform 1 0 552 0 1 1079
box -32 -26 32 26
use via_M3_M4_0  NoName_53
timestamp 1704387757
transform 1 0 276 0 1 1079
box -32 -26 32 26
use via_M3_M4_0  NoName_55
timestamp 1704387757
transform 1 0 1656 0 1 1079
box -32 -26 32 26
use via_M3_M4_0  NoName_57
timestamp 1704387757
transform 1 0 1932 0 1 1079
box -32 -26 32 26
use via_M4_M5_0  NoName_60
timestamp 1706182685
transform 1 0 2576 0 1 1162
box -37 -34 37 34
use via_M4_M5_0  NoName_62
timestamp 1706182685
transform 1 0 2576 0 1 415
box -37 -34 37 34
use via_M3_M4_0  NoName_64
timestamp 1704387757
transform 1 0 2760 0 1 1162
box -32 -26 32 26
use via_M3_M4_0  NoName_65
timestamp 1704387757
transform 1 0 6440 0 1 415
box -32 -26 32 26
use via_M3_M4_0  NoName_66
timestamp 1704387757
transform 1 0 5980 0 1 1328
box -32 -26 32 26
use via_M3_M4_0  NoName_68
timestamp 1704387757
transform 1 0 7176 0 1 1328
box -32 -26 32 26
use via_M3_M4_0  NoName_70
timestamp 1704387757
transform 1 0 6072 0 1 1328
box -32 -26 32 26
use via_M3_M4_0  NoName_72
timestamp 1704387757
transform 1 0 7360 0 1 1328
box -32 -26 32 26
use via_M3_M4_0  NoName_76
timestamp 1704387757
transform 1 0 7912 0 1 1162
box -32 -26 32 26
use via_M3_M4_0  NoName_78
timestamp 1704387757
transform 1 0 8280 0 1 996
box -32 -26 32 26
use via_M4_M5_0  NoName_81
timestamp 1706182685
transform 1 0 8096 0 1 996
box -37 -34 37 34
use via_M4_M5_0  NoName_83
timestamp 1706182685
transform 1 0 8096 0 1 581
box -37 -34 37 34
use via_M3_M4_0  NoName_85
timestamp 1704387757
transform 1 0 8372 0 1 581
box -32 -26 32 26
use via_M3_M4_0  NoName_88
timestamp 1704387757
transform 1 0 8280 0 1 498
box -32 -26 32 26
use via_M3_M4_0  NoName_90
timestamp 1704387757
transform 1 0 8556 0 1 498
box -32 -26 32 26
use via_M3_M4_0  NoName_93
timestamp 1704387757
transform 1 0 8832 0 1 581
box -32 -26 32 26
use via_M3_M4_0  NoName_95
timestamp 1704387757
transform 1 0 9108 0 1 581
box -32 -26 32 26
use via_M4_M5_0  NoName_98
timestamp 1706182685
transform 1 0 9568 0 1 581
box -37 -34 37 34
use via_M4_M5_0  NoName_100
timestamp 1706182685
transform 1 0 9568 0 1 1162
box -37 -34 37 34
use via_M3_M4_0  NoName_102
timestamp 1704387757
transform 1 0 9752 0 1 581
box -32 -26 32 26
use via_M3_M4_0  NoName_103
timestamp 1704387757
transform 1 0 10028 0 1 1162
box -32 -26 32 26
use via_M3_M4_0  via_M3_M4_0_0
timestamp 1704387757
transform 1 0 5704 0 1 1162
box -32 -26 32 26
<< labels >>
flabel metal1 1380 1245 1380 1245 0 FreeSans 512 90 0 0 SCAN_CLK
port 1 nsew
flabel metal1 184 1245 184 1245 0 FreeSans 512 90 0 0 SCAN_CLK_OUT
port 2 nsew
flabel metal1 2024 415 2024 415 0 FreeSans 512 90 0 0 SCAN_DATA_IN
port 3 nsew
flabel metal1 8648 1245 8648 1245 0 FreeSans 512 90 0 0 SCAN_DATA_OUT
port 4 nsew
flabel metal1 1564 1245 1564 1245 0 FreeSans 512 90 0 0 SCAN_EN
port 5 nsew
flabel metal1 7176 1245 7176 1245 0 FreeSans 512 90 0 0 SCAN_GATE
port 6 nsew
flabel metal1 6440 1245 6440 1245 0 FreeSans 512 90 0 0 SCAN_GATE_VALUE
port 7 nsew
flabel metal1 552 415 552 415 0 FreeSans 512 90 0 0 SCAN_IN
port 8 nsew
flabel metal1 92 415 92 415 0 FreeSans 512 90 0 0 SCAN_LOAD
port 9 nsew
flabel metal1 7912 415 7912 415 0 FreeSans 512 90 0 0 SCAN_OUT
port 10 nsew
<< end >>
