magic
tech sky130A
magscale 1 2
timestamp 1646748542
<< nwell >>
rect -66 208 234 448
<< pmos >>
rect 29 244 59 412
rect 115 244 145 412
<< pdiff >>
rect -24 381 29 412
rect -24 347 -16 381
rect 18 347 29 381
rect -24 309 29 347
rect -24 275 -16 309
rect 18 275 29 309
rect -24 244 29 275
rect 59 381 115 412
rect 59 347 70 381
rect 104 347 115 381
rect 59 309 115 347
rect 59 275 70 309
rect 104 275 115 309
rect 59 244 115 275
rect 145 381 198 412
rect 145 347 156 381
rect 190 347 198 381
rect 145 309 198 347
rect 145 275 156 309
rect 190 275 198 309
rect 145 244 198 275
<< pdiffc >>
rect -16 347 18 381
rect -16 275 18 309
rect 70 347 104 381
rect 70 275 104 309
rect 156 347 190 381
rect 156 275 190 309
<< poly >>
rect 20 495 154 511
rect 20 461 36 495
rect 70 461 104 495
rect 138 461 154 495
rect 20 443 154 461
rect 29 438 145 443
rect 29 412 59 438
rect 115 412 145 438
rect 29 218 59 244
rect 115 218 145 244
< polycont >>
rect 36 461 70 495
rect 104 461 138 495
<< locali >>
rect 20 495 154 511
rect 20 461 34 495
rect 70 461 104 495
rect 140 461 154 495
rect 20 443 154 461
rect -16 381 18 397
rect -16 309 18 347
rect -16 259 18 275
rect 70 381 104 397
rect 70 309 104 347
rect 70 259 104 275
rect 156 381 190 397
rect 156 309 190 347
rect 156 259 190 275
<< viali >>
rect 34 461 36 495
rect 36 461 68 495
rect 106 461 138 495
rect 138 461 140 495
rect -16 347 18 381
rect -16 275 18 309
rect 70 347 104 381
rect 70 275 104 309
rect 156 347 190 381
rect 156 275 190 309
<< metal1 >>
rect 22 495 152 507
rect 22 461 34 495
rect 68 461 106 495
rect 140 461 152 495
rect 22 449 152 461
rect -22 381 24 397
rect -22 347 -16 381
rect 18 347 24 381
rect -22 309 24 347
rect -22 275 -16 309
rect 18 275 24 309
rect -22 179 24 275
rect 61 386 113 397
rect 61 322 113 334
rect 61 259 113 270
rect 150 381 196 397
rect 150 347 156 381
rect 190 347 196 381
rect 150 309 196 347
rect 150 275 156 309
rect 190 275 196 309
rect 150 179 196 275
rect -22 119 196 179
<< via1 >>
rect 61 381 113 386
rect 61 347 70 381
rect 70 347 104 381
rect 104 347 113 381
rect 61 334 113 347
rect 61 309 113 322
rect 61 275 70 309
rect 70 275 104 309
rect 104 275 113 309
rect 61 270 113 275
<< metal2 >>
rect 61 386 113 392
rect 61 322 113 334
rect 61 264 113 270
<< end >>
