magic
tech sky130A
magscale 1 2
timestamp 1679560816
<< checkpaint >>
rect -1300 -1325 3604 3337
<< metal1 >>
rect 114 1688 174 2056
rect 402 1688 462 2056
rect 690 1688 750 2056
rect 978 1688 1038 2056
rect 1266 1688 1326 2056
rect 1554 1688 1614 2056
rect 1842 1688 1902 2056
rect 2130 1688 2190 2056
rect 114 -40 174 328
rect 402 -40 462 328
rect 690 -40 750 328
rect 978 -40 1038 328
rect 1266 -40 1326 328
rect 1554 -40 1614 328
rect 1842 -40 1902 328
rect 2130 -40 2190 328
<< metal2 >>
rect -40 1956 2344 2076
rect 212 1554 2092 1614
rect 124 1266 2092 1326
rect 124 690 2092 750
rect 212 402 2092 462
rect -40 -60 2344 60
<< metal3 >>
rect 114 690 174 1326
rect 258 432 318 1584
rect 546 432 606 1584
rect 834 432 894 1584
rect 1122 432 1182 1584
rect 1410 432 1470 1584
rect 1698 432 1758 1584
rect 1986 402 2046 1614
use nmos13_fast_boundary  MN0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 144 1008
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 2160 0 1 0
box 0 0 144 1008
use nmos13_fast_center_nf2  MN0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 6 288 0 0 1008
timestamp 1654175211
transform 1 0 144 0 1 0
box -92 286 380 756
use via_M1_M2_0  MN0_IVD0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 6 288 0 0 1008
timestamp 1647525606
transform 1 0 288 0 1 432
box -32 -32 32 32
use via_M1_M2_0  MN0_IVG0
array 0 6 288 0 0 1008
timestamp 1647525606
transform 1 0 288 0 1 720
box -32 -32 32 32
use via_M1_M2_1  MN0_IVTIED0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 7 288 0 0 1008
timestamp 1647525606
transform 1 0 144 0 1 0
box -32 -32 32 32
use pmos13_fast_boundary  MP0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 2016
box 0 0 144 1008
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 2160 0 -1 2016
box 0 0 144 1008
use pmos13_fast_center_nf2  MP0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 6 288 0 0 -1008
timestamp 1654091791
transform 1 0 144 0 -1 2016
box -92 132 380 756
use via_M1_M2_0  MP0_IVD0
array 0 6 288 0 0 -1008
timestamp 1647525606
transform 1 0 288 0 -1 1584
box -32 -32 32 32
use via_M1_M2_0  MP0_IVG0
array 0 6 288 0 0 -1008
timestamp 1647525606
transform 1 0 288 0 -1 1296
box -32 -32 32 32
use via_M1_M2_1  MP0_IVTIED0
array 0 7 288 0 0 -1008
timestamp 1647525606
transform 1 0 144 0 -1 2016
box -32 -32 32 32
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 144 0 1 720
box -38 -38 38 38
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 144 0 1 1296
box -38 -38 38 38
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 2016 0 1 432
box -38 -38 38 38
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 2016 0 1 1584
box -38 -38 38 38
<< labels >>
flabel metal3 144 1008 144 1008 0 FreeSans 480 90 0 0 I
port 7 nsew
flabel metal3 288 1008 288 1008 0 FreeSans 480 90 0 0 O
port 8 nsew
flabel metal3 576 1008 576 1008 0 FreeSans 480 90 0 0 O
port 9 nsew
flabel metal3 864 1008 864 1008 0 FreeSans 480 90 0 0 O
port 10 nsew
flabel metal3 1152 1008 1152 1008 0 FreeSans 480 90 0 0 O
port 11 nsew
flabel metal3 1440 1008 1440 1008 0 FreeSans 480 90 0 0 O
port 12 nsew
flabel metal3 1728 1008 1728 1008 0 FreeSans 480 90 0 0 O
port 13 nsew
flabel metal3 2016 1008 2016 1008 0 FreeSans 480 90 0 0 O
port 14 nsew
flabel metal2 288 2016 288 2016 0 FreeSans 960 0 0 0 VDD
port 15 nsew
flabel metal2 432 2016 432 2016 0 FreeSans 960 0 0 0 VDD
port 16 nsew
flabel metal2 576 2016 576 2016 0 FreeSans 960 0 0 0 VDD
port 17 nsew
flabel metal2 720 2016 720 2016 0 FreeSans 960 0 0 0 VDD
port 18 nsew
flabel metal2 864 2016 864 2016 0 FreeSans 960 0 0 0 VDD
port 19 nsew
flabel metal2 1008 2016 1008 2016 0 FreeSans 960 0 0 0 VDD
port 20 nsew
flabel metal2 1152 2016 1152 2016 0 FreeSans 960 0 0 0 VDD
port 21 nsew
flabel metal2 288 0 288 0 0 FreeSans 960 0 0 0 VSS
port 22 nsew
flabel metal2 432 0 432 0 0 FreeSans 960 0 0 0 VSS
port 23 nsew
flabel metal2 576 0 576 0 0 FreeSans 960 0 0 0 VSS
port 24 nsew
flabel metal2 720 0 720 0 0 FreeSans 960 0 0 0 VSS
port 25 nsew
flabel metal2 864 0 864 0 0 FreeSans 960 0 0 0 VSS
port 26 nsew
flabel metal2 1008 0 1008 0 0 FreeSans 960 0 0 0 VSS
port 27 nsew
flabel metal2 1152 0 1152 0 0 FreeSans 960 0 0 0 VSS
port 28 nsew
<< end >>
