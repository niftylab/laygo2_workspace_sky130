** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/dec_3to8.sch
.subckt dec_3to8 A2 A1 A0 VDD VSS O0 O1 O2 O3 O4 O5 O6 O7 EN
*.PININFO A2:I A1:I A0:I VDD:B VSS:B O0:O O1:O O2:O O3:O O4:O O5:O O6:O O7:O EN:I
X_inv7 A2 VDD VSS net3 inv NF=2
X_inv1 A1 VDD VSS net2 inv NF=2
X_inv2 A0 VDD VSS net1 inv NF=2
x_AndF1 net3 net2 O0 VDD VSS net1 EN and_4in NF=2
x_AndF2 net3 net2 O1 VDD VSS A0 EN and_4in NF=2
x_AndF7 A2 A1 O6 VDD VSS net1 EN and_4in NF=2
x_AndF8 A2 A1 O7 VDD VSS A0 EN and_4in NF=2
x_AndF3 net3 A1 O2 VDD VSS net1 EN and_4in NF=2
x_AndF4 net3 A1 O3 VDD VSS A0 EN and_4in NF=2
x_AndF5 A2 net2 O4 VDD VSS net1 EN and_4in NF=2
x_AndF6 A2 net2 O5 VDD VSS A0 EN and_4in NF=2
.ends

* expanding   symbol:
*+  /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/inv.sym # of pins=4
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/inv.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/inv.sch
.subckt inv X VDD VSS Y  NF=2
*.PININFO VSS:B X:I Y:O VDD:B
XM1 Y X VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM2 Y X VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
.ends


* expanding   symbol:
*+  /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/and_4in.sym # of pins=7
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/and_4in.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/and_4in.sch
.subckt and_4in B D O VDD VSS C A  NF=2
*.PININFO VDD:B VSS:B A:I B:I C:I D:I O:O
X_nand2 D C net2 VDD VSS nand NF=2
X_nand1 B A net1 VDD VSS nand NF=2
X_nand3 O net1 net2 VDD VSS nor NF=2
.ends


* expanding   symbol:
*+  /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nand.sym # of pins=5
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nand.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nand.sch
.subckt nand B A Y VDD VSS  NF=2
*.PININFO Y:O A:I VDD:B VSS:B B:I
XM1 Y A net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM2 net1 B VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM3 Y B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
XM4 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
.ends


* expanding   symbol:
*+  /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nor.sym # of pins=5
** sym_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nor.sym
** sch_path:
*+ /Users/brianlsy/Desktop/brianlsy/git_workspace/fork/laygo2_workspace_sky130/xschem_lib/sylee21/nor.sch
.subckt nor Y A B VDD VSS  NF=2
*.PININFO VDD:B VSS:B Y:O A:I B:I
XM1 Y B VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1 m=NF
XM3 Y A net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
XM4 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=1 m=NF
.ends

.end
