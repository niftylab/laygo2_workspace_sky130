magic
tech sky130A
magscale 1 2
timestamp 1706249518
<< checkpaint >>
rect -1260 2124 2072 2156
rect -1294 -799 2072 2124
rect -1294 -1294 2030 -799
rect -1260 -1344 1996 -1294
<< locali >>
rect 66 730 118 847
rect 250 730 302 847
rect 342 730 689 764
rect 342 598 394 730
rect 150 564 394 598
rect 518 564 586 598
rect 150 481 218 515
rect 443 481 586 515
rect 150 315 218 349
rect 518 315 661 349
rect 150 232 394 266
rect 518 232 586 266
rect 342 100 394 232
rect 66 -17 118 100
rect 250 -17 302 100
rect 342 66 689 100
<< metal1 >>
rect -17 804 753 856
rect 152 306 216 524
rect 428 306 492 524
rect 520 223 584 607
rect 612 306 676 524
rect -17 -26 753 26
use nmos130_fast_boundary  MN0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363493
transform 1 0 0 0 1 0
box 0 -84 92 280
use nmos130_fast_boundary  MN0_IBNDR0
timestamp 1704363493
transform 1 0 276 0 1 0
box 0 -84 92 280
use nmos130_fast_center_nf2  MN0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704390143
transform 1 0 92 0 1 0
box -31 -84 215 362
use via_M1_M2_0  MN0_IVD0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704392934
transform 1 0 184 0 1 249
box -17 -17 17 17
use via_M1_M2_0  MN0_IVG0
timestamp 1704392934
transform 1 0 184 0 1 332
box -17 -17 17 17
use via_M1_M2_1  MN0_IVTIED0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 184 0 0 415
timestamp 1704386328
transform 1 0 92 0 1 0
box -26 -26 26 26
use nmos130_fast_boundary  MN1_IBNDL0
timestamp 1704363493
transform 1 0 368 0 1 0
box 0 -84 92 280
use nmos130_fast_boundary  MN1_IBNDR0
timestamp 1704363493
transform 1 0 644 0 1 0
box 0 -84 92 280
use nmos130_fast_center_nf2  MN1_IM0
timestamp 1704390143
transform 1 0 460 0 1 0
box -31 -84 215 362
use via_M1_M2_0  MN1_IVD0
timestamp 1704392934
transform 1 0 552 0 1 249
box -17 -17 17 17
use via_M1_M2_0  MN1_IVG0
timestamp 1704392934
transform 1 0 552 0 1 332
box -17 -17 17 17
use via_M1_M2_0  MN1_IVS0
array 0 1 184 0 0 415
timestamp 1704392934
transform 1 0 460 0 1 83
box -17 -17 17 17
use pmos130_fast_boundary  MP0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363574
transform 1 0 0 0 -1 830
box 0 -66 168 369
use pmos130_fast_boundary  MP0_IBNDR0
timestamp 1704363574
transform 1 0 276 0 -1 830
box 0 -66 168 369
use pmos130_fast_center_nf2  MP0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704364343
transform 1 0 92 0 -1 830
box -31 -66 215 369
use via_M1_M2_0  MP0_IVD0
timestamp 1704392934
transform 1 0 184 0 -1 581
box -17 -17 17 17
use via_M1_M2_0  MP0_IVG0
timestamp 1704392934
transform 1 0 184 0 -1 498
box -17 -17 17 17
use via_M1_M2_1  MP0_IVTIED0
array 0 1 184 0 0 -415
timestamp 1704386328
transform 1 0 92 0 -1 830
box -26 -26 26 26
use pmos130_fast_boundary  MP1_IBNDL0
timestamp 1704363574
transform 1 0 368 0 -1 830
box 0 -66 168 369
use pmos130_fast_boundary  MP1_IBNDR0
timestamp 1704363574
transform 1 0 644 0 -1 830
box 0 -66 168 369
use pmos130_fast_center_nf2  MP1_IM0
timestamp 1704364343
transform 1 0 460 0 -1 830
box -31 -66 215 369
use via_M1_M2_0  MP1_IVD0
timestamp 1704392934
transform 1 0 552 0 -1 581
box -17 -17 17 17
use via_M1_M2_0  MP1_IVG0
timestamp 1704392934
transform 1 0 552 0 -1 498
box -17 -17 17 17
use via_M1_M2_0  MP1_IVS0
array 0 1 184 0 0 -415
timestamp 1704392934
transform 1 0 460 0 -1 747
box -17 -17 17 17
use via_M2_M3_0  NoName_0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704386899
transform 1 0 184 0 1 332
box -32 -17 32 17
use via_M2_M3_0  NoName_2
timestamp 1704386899
transform 1 0 184 0 1 498
box -32 -17 32 17
use via_M2_M3_0  NoName_3
timestamp 1704386899
transform 1 0 552 0 1 249
box -32 -17 32 17
use via_M2_M3_0  NoName_5
timestamp 1704386899
transform 1 0 552 0 1 581
box -32 -17 32 17
use via_M2_M3_0  NoName_6
timestamp 1704386899
transform 1 0 644 0 1 332
box -32 -17 32 17
use via_M2_M3_0  NoName_10
timestamp 1704386899
transform 1 0 460 0 1 498
box -32 -17 32 17
use via_M1_M2_0  NoName_13
timestamp 1704392934
transform 1 0 368 0 1 581
box -17 -17 17 17
use via_M1_M2_0  NoName_15
timestamp 1704392934
transform 1 0 368 0 1 747
box -17 -17 17 17
use via_M1_M2_0  NoName_18
timestamp 1704392934
transform 1 0 368 0 1 249
box -17 -17 17 17
use via_M1_M2_0  NoName_20
timestamp 1704392934
transform 1 0 368 0 1 83
box -17 -17 17 17
<< labels >>
flabel metal1 644 415 644 415 0 FreeSans 512 90 0 0 EN
port 1 nsew
flabel metal1 460 415 460 415 0 FreeSans 512 90 0 0 ENB
port 2 nsew
flabel metal1 184 415 184 415 0 FreeSans 512 90 0 0 I
port 3 nsew
flabel metal1 552 415 552 415 0 FreeSans 512 90 0 0 O
port 4 nsew
flabel metal1 368 830 368 830 0 FreeSans 416 0 0 0 VDD
port 5 nsew
flabel metal1 368 0 368 0 0 FreeSans 416 0 0 0 VSS
port 6 nsew
<< end >>
