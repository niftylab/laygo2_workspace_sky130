magic
tech sky130A
timestamp 1654176175
<< nwell >>
rect -46 66 190 342
<< pmos >>
rect 28 84 43 324
rect 100 84 115 324
<< pdiff >>
rect -28 289 28 324
rect -28 269 -10 289
rect 10 269 28 289
rect -28 239 28 269
rect -28 219 -10 239
rect 10 219 28 239
rect -28 189 28 219
rect -28 169 -10 189
rect 10 169 28 189
rect -28 139 28 169
rect -28 119 -10 139
rect 10 119 28 139
rect -28 84 28 119
rect 43 289 100 324
rect 43 269 62 289
rect 82 269 100 289
rect 43 239 100 269
rect 43 219 62 239
rect 82 219 100 239
rect 43 189 100 219
rect 43 169 62 189
rect 82 169 100 189
rect 43 139 100 169
rect 43 119 62 139
rect 82 119 100 139
rect 43 84 100 119
rect 115 289 172 324
rect 115 269 134 289
rect 154 269 172 289
rect 115 239 172 269
rect 115 219 134 239
rect 154 219 172 239
rect 115 189 172 219
rect 115 169 134 189
rect 154 169 172 189
rect 115 139 172 169
rect 115 119 134 139
rect 154 119 172 139
rect 115 84 172 119
<< pdiffc >>
rect -10 269 10 289
rect -10 219 10 239
rect -10 169 10 189
rect -10 119 10 139
rect 62 269 82 289
rect 62 219 82 239
rect 62 169 82 189
rect 62 119 82 139
rect 134 269 154 289
rect 134 219 154 239
rect 134 169 154 189
rect 134 119 154 139
<< poly >>
rect -17 369 43 378
rect -17 351 -6 369
rect 12 351 43 369
rect -17 342 43 351
rect 28 324 43 342
rect 100 369 160 378
rect 100 351 136 369
rect 154 351 160 369
rect 100 342 160 351
rect 100 324 115 342
rect 28 66 43 84
rect 100 66 115 84
<< polycont >>
rect -6 351 12 369
rect 136 351 154 369
<< locali >>
rect -17 369 28 378
rect -17 351 -6 369
rect 12 351 28 369
rect -17 342 28 351
rect 115 369 160 378
rect 115 351 136 369
rect 154 351 160 369
rect 115 342 160 351
rect -15 289 15 297
rect -15 269 -10 289
rect 10 269 15 289
rect -15 239 15 269
rect -15 219 -10 239
rect 10 219 15 239
rect -15 189 15 219
rect -15 169 -10 189
rect 10 169 15 189
rect -15 139 15 169
rect -15 119 -10 139
rect 10 119 15 139
rect -15 111 15 119
rect 57 289 87 297
rect 57 269 62 289
rect 82 269 87 289
rect 57 239 87 269
rect 57 219 62 239
rect 82 219 87 239
rect 57 189 87 219
rect 57 169 62 189
rect 82 169 87 189
rect 57 139 87 169
rect 57 119 62 139
rect 82 119 87 139
rect 57 111 87 119
rect 129 289 159 297
rect 129 269 134 289
rect 154 269 159 289
rect 129 239 159 269
rect 129 219 134 239
rect 154 219 159 239
rect 129 189 159 219
rect 129 169 134 189
rect 154 169 159 189
rect 129 139 159 169
rect 129 119 134 139
rect 154 119 159 139
rect 129 111 159 119
<< viali >>
rect -6 351 12 369
rect 136 351 154 369
rect -10 269 10 289
rect -10 219 10 239
rect -10 169 10 189
rect -10 119 10 139
rect 62 269 82 289
rect 62 219 82 239
rect 62 169 82 189
rect 62 119 82 139
rect 134 269 154 289
rect 134 219 154 239
rect 134 169 154 189
rect 134 119 154 139
<< metal1 >>
rect -17 369 28 378
rect -17 351 -6 369
rect 12 351 28 369
rect -17 342 28 351
rect 115 369 160 378
rect 115 351 136 369
rect 154 351 160 369
rect 115 342 160 351
rect -15 289 15 297
rect -15 269 -10 289
rect 10 269 15 289
rect -15 239 15 269
rect -15 219 -10 239
rect 10 219 15 239
rect -15 189 15 219
rect -15 169 -10 189
rect 10 169 15 189
rect -15 139 15 169
rect -15 119 -10 139
rect 10 119 15 139
rect -15 94 15 119
rect 57 289 87 297
rect 57 269 62 289
rect 82 269 87 289
rect 57 239 87 269
rect 57 219 62 239
rect 82 219 87 239
rect 57 189 87 219
rect 57 169 62 189
rect 82 169 87 189
rect 57 139 87 169
rect 57 119 62 139
rect 82 119 87 139
rect 57 94 87 119
rect 129 289 159 297
rect 129 269 134 289
rect 154 269 159 289
rect 129 239 159 269
rect 129 219 134 239
rect 154 219 159 239
rect 129 189 159 219
rect 129 169 134 189
rect 154 169 159 189
rect 129 139 159 169
rect 129 119 134 139
rect 154 119 159 139
rect 129 94 159 119
<< labels >>
flabel metal1 -17 342 28 378 0 FreeSans 80 0 0 0 G0
port 2 nsew
flabel metal1 115 342 160 378 0 FreeSans 80 0 0 0 G1
port 3 nsew
flabel metal1 -15 94 15 297 0 FreeSans 80 0 0 0 S0
port 4 nsew
flabel nwell -10 327 2 335 0 FreeSans 40 0 0 0 BODY
port 6 nsew
flabel metal1 129 94 159 297 0 FreeSans 80 0 0 0 D0
port 1 e
<< end >>
