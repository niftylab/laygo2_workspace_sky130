magic
tech sky130A
timestamp 1679561058
<< checkpaint >>
rect -650 -660 2378 1668
<< metal2 >>
rect -20 978 1748 1038
rect 993 129 1527 159
rect 417 57 1311 87
rect -20 -30 1748 30
<< metal3 >>
rect 129 360 159 648
rect 345 360 375 648
rect 705 360 735 648
rect 921 360 951 648
rect 417 57 447 159
rect 1281 57 1311 375
rect 1497 129 1527 375
rect 1569 216 1599 864
use logic_generated_nand_2x  nand0 magic_layout/logic_generated
timestamp 1679560872
transform 1 0 0 0 1 0
box -20 -30 596 1038
use logic_generated_nand_2x  nand1
timestamp 1679560872
transform 1 0 576 0 1 0
box -20 -30 596 1038
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 432 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 1296 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 1008 0 1 144
box -19 -19 19 19
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 1512 0 1 144
box -19 -19 19 19
use logic_generated_nor_2x  nor0 magic_layout/logic_generated
timestamp 1679560883
transform 1 0 1152 0 1 0
box -20 -30 596 1038
<< labels >>
flabel metal3 936 504 936 504 0 FreeSans 240 90 0 0 A
port 1 nsew
flabel metal3 720 504 720 504 0 FreeSans 240 90 0 0 B
port 2 nsew
flabel metal3 360 504 360 504 0 FreeSans 240 90 0 0 C
port 3 nsew
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 D
port 4 nsew
flabel metal2 864 1008 864 1008 0 FreeSans 480 0 0 0 VDD
port 5 nsew
flabel metal2 864 0 864 0 0 FreeSans 480 0 0 0 VSS
port 6 nsew
flabel metal3 1584 540 1584 540 0 FreeSans 240 90 0 0 Y
port 7 nsew
<< end >>
