magic
tech sky130A
timestamp 1679560843
<< checkpaint >>
rect -650 -660 1514 1668
<< metal2 >>
rect -20 978 884 1038
rect 273 489 519 519
rect -20 -30 884 30
<< metal3 >>
rect 57 360 87 648
rect 273 201 303 519
rect 489 345 519 519
rect 705 216 735 792
use logic_generated_inv_4x  inv0 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 0 0 1 0
box -20 -30 452 1038
use logic_generated_inv_4x  inv1
timestamp 1679560816
transform 1 0 432 0 1 0
box -20 -30 452 1038
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 288 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 504 0 1 504
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 I
port 1 nsew
flabel metal3 720 504 720 504 0 FreeSans 240 90 0 0 O
port 2 nsew
flabel metal2 432 1008 432 1008 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal2 432 0 432 0 0 FreeSans 480 0 0 0 VSS
port 4 nsew
<< end >>
