magic
tech sky130A
timestamp 1679561070
<< checkpaint >>
rect -650 -660 5834 1668
<< metal2 >>
rect -20 978 5204 1038
rect 129 849 2175 879
rect 57 489 4479 519
rect 345 417 4695 447
rect 1281 273 1527 303
rect 2433 273 2679 303
rect 3585 273 3831 303
rect 4737 273 4983 303
rect 417 57 3543 87
rect -20 -30 5204 30
<< metal3 >>
rect 57 345 87 648
rect 129 216 159 879
rect 345 345 375 648
rect 417 57 447 792
rect 993 633 1023 879
rect 1209 57 1239 375
rect 1281 201 1311 303
rect 1497 273 1527 375
rect 1569 216 1599 792
rect 2145 633 2175 879
rect 2361 345 2391 447
rect 2433 201 2463 303
rect 2649 273 2679 375
rect 2721 216 2751 792
rect 3297 345 3327 519
rect 3513 57 3543 375
rect 3585 201 3615 303
rect 3801 273 3831 375
rect 3873 216 3903 792
rect 4449 345 4479 519
rect 4665 345 4695 447
rect 4737 201 4767 303
rect 4953 273 4983 375
rect 5025 216 5055 792
<< metal4 >>
rect 705 345 4191 375
use logic_generated_inv_2x  inv0 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 0 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv1
timestamp 1679560816
transform 1 0 288 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv_0
timestamp 1679560816
transform 1 0 1440 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv_1
timestamp 1679560816
transform 1 0 2592 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv_2
timestamp 1679560816
transform 1 0 3744 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv_3
timestamp 1679560816
transform 1 0 4896 0 1 0
box -20 -30 308 1038
use logic_generated_nand3_2x  nand3_0 magic_layout/logic_generated
timestamp 1679560960
transform 1 0 576 0 1 0
box -20 -30 884 1038
use logic_generated_nand3_2x  nand3_1
timestamp 1679560960
transform 1 0 1728 0 1 0
box -20 -30 884 1038
use logic_generated_nand3_2x  nand3_2
timestamp 1679560960
transform 1 0 2880 0 1 0
box -20 -30 884 1038
use logic_generated_nand3_2x  nand3_3
timestamp 1679560960
transform 1 0 4032 0 1 0
box -20 -30 884 1038
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 432 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 1224 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 3528 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_8
timestamp 1647525786
transform 1 0 360 0 1 432
box -19 -19 19 19
use via_M2_M3_0  NoName_10
timestamp 1647525786
transform 1 0 2376 0 1 432
box -19 -19 19 19
use via_M2_M3_0  NoName_12
timestamp 1647525786
transform 1 0 4680 0 1 432
box -19 -19 19 19
use via_M2_M3_0  NoName_15
timestamp 1647525786
transform 1 0 144 0 1 864
box -19 -19 19 19
use via_M2_M3_0  NoName_17
timestamp 1647525786
transform 1 0 1008 0 1 864
box -19 -19 19 19
use via_M2_M3_0  NoName_19
timestamp 1647525786
transform 1 0 2160 0 1 864
box -19 -19 19 19
use via_M2_M3_0  NoName_22
timestamp 1647525786
transform 1 0 72 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_24
timestamp 1647525786
transform 1 0 3312 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_26
timestamp 1647525786
transform 1 0 4464 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_29
timestamp 1647525786
transform 1 0 1296 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_31
timestamp 1647525786
transform 1 0 1512 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_34
timestamp 1647525786
transform 1 0 2448 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_36
timestamp 1647525786
transform 1 0 2664 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_39
timestamp 1647525786
transform 1 0 3600 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_41
timestamp 1647525786
transform 1 0 3816 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_44
timestamp 1647525786
transform 1 0 4752 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_46
timestamp 1647525786
transform 1 0 4968 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_48 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 720 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_49
timestamp 1647526059
transform 1 0 1872 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_50
timestamp 1647526059
transform 1 0 3024 0 1 360
box -19 -19 19 19
use via_M3_M4_0  NoName_51
timestamp 1647526059
transform 1 0 4176 0 1 360
box -19 -19 19 19
<< labels >>
flabel metal3 360 504 360 504 0 FreeSans 240 90 0 0 A0
port 1 nsew
flabel metal3 432 504 432 504 0 FreeSans 240 90 0 0 A0bar
port 2 nsew
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 A1
port 3 nsew
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 A1bar
port 4 nsew
flabel metal4 2448 360 2448 360 0 FreeSans 240 0 0 0 EN
port 5 nsew
flabel metal2 2592 1008 2592 1008 0 FreeSans 480 0 0 0 VDD
port 6 nsew
flabel metal2 2592 0 2592 0 0 FreeSans 480 0 0 0 VSS
port 7 nsew
flabel metal3 1584 504 1584 504 0 FreeSans 240 90 0 0 Y0
port 8 nsew
flabel metal3 2736 504 2736 504 0 FreeSans 240 90 0 0 Y1
port 9 nsew
flabel metal3 3888 504 3888 504 0 FreeSans 240 90 0 0 Y2
port 10 nsew
flabel metal3 5040 504 5040 504 0 FreeSans 240 90 0 0 Y3
port 11 nsew
<< end >>
