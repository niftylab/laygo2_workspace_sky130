magic
tech sky130A
magscale 1 2
timestamp 1706178735
<< checkpaint >>
rect -1260 2124 2440 2156
rect -1294 -799 2440 2124
rect -1294 -1294 2398 -799
rect -1260 -1344 2364 -1294
<< locali >>
rect 66 713 118 864
rect 250 713 302 864
rect 434 713 486 864
rect 526 730 1057 764
rect 526 598 578 730
rect 139 564 578 598
rect 691 564 965 598
rect 139 481 413 515
rect 691 481 965 515
rect 139 315 413 349
rect 691 315 1029 349
rect 139 232 578 266
rect 691 232 965 266
rect 66 -34 118 117
rect 250 -34 302 117
rect 434 -34 486 117
rect 526 100 578 232
rect 526 66 1057 100
<< metal1 >>
rect -34 804 1138 856
rect 152 306 216 524
rect 796 306 860 524
rect 888 223 952 607
rect 980 306 1044 524
rect -34 -26 1138 26
use nmos130_fast_boundary  MN0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363493
transform 1 0 0 0 1 0
box 0 -84 92 280
use nmos130_fast_boundary  MN0_IBNDR0
timestamp 1704363493
transform 1 0 460 0 1 0
box 0 -84 92 280
use nmos130_fast_center_nf2  MN0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 184 0 0 415
timestamp 1704390143
transform 1 0 92 0 1 0
box -31 -84 215 362
use via_M1_M2_0  MN0_IVD0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 184 0 0 415
timestamp 1704392934
transform 1 0 184 0 1 249
box -17 -17 17 17
use via_M1_M2_0  MN0_IVG0
array 0 1 184 0 0 415
timestamp 1704392934
transform 1 0 184 0 1 332
box -17 -17 17 17
use via_M1_M2_1  MN0_IVTIED0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 2 184 0 0 415
timestamp 1704386328
transform 1 0 92 0 1 0
box -26 -26 26 26
use nmos130_fast_boundary  MN1_IBNDL0
timestamp 1704363493
transform 1 0 552 0 1 0
box 0 -84 92 280
use nmos130_fast_boundary  MN1_IBNDR0
timestamp 1704363493
transform 1 0 1012 0 1 0
box 0 -84 92 280
use nmos130_fast_center_nf2  MN1_IM0
array 0 1 184 0 0 415
timestamp 1704390143
transform 1 0 644 0 1 0
box -31 -84 215 362
use via_M1_M2_0  MN1_IVD0
array 0 1 184 0 0 415
timestamp 1704392934
transform 1 0 736 0 1 249
box -17 -17 17 17
use via_M1_M2_0  MN1_IVG0
array 0 1 184 0 0 415
timestamp 1704392934
transform 1 0 736 0 1 332
box -17 -17 17 17
use via_M1_M2_0  MN1_IVS0
array 0 2 184 0 0 415
timestamp 1704392934
transform 1 0 644 0 1 83
box -17 -17 17 17
use pmos130_fast_boundary  MP0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363574
transform 1 0 0 0 -1 830
box 0 -66 168 369
use pmos130_fast_boundary  MP0_IBNDR0
timestamp 1704363574
transform 1 0 460 0 -1 830
box 0 -66 168 369
use pmos130_fast_center_nf2  MP0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 184 0 0 -415
timestamp 1704364343
transform 1 0 92 0 -1 830
box -31 -66 215 369
use via_M1_M2_0  MP0_IVD0
array 0 1 184 0 0 -415
timestamp 1704392934
transform 1 0 184 0 -1 581
box -17 -17 17 17
use via_M1_M2_0  MP0_IVG0
array 0 1 184 0 0 -415
timestamp 1704392934
transform 1 0 184 0 -1 498
box -17 -17 17 17
use via_M1_M2_1  MP0_IVTIED0
array 0 2 184 0 0 -415
timestamp 1704386328
transform 1 0 92 0 -1 830
box -26 -26 26 26
use pmos130_fast_boundary  MP1_IBNDL0
timestamp 1704363574
transform 1 0 552 0 -1 830
box 0 -66 168 369
use pmos130_fast_boundary  MP1_IBNDR0
timestamp 1704363574
transform 1 0 1012 0 -1 830
box 0 -66 168 369
use pmos130_fast_center_nf2  MP1_IM0
array 0 1 184 0 0 -415
timestamp 1704364343
transform 1 0 644 0 -1 830
box -31 -66 215 369
use via_M1_M2_0  MP1_IVD0
array 0 1 184 0 0 -415
timestamp 1704392934
transform 1 0 736 0 -1 581
box -17 -17 17 17
use via_M1_M2_0  MP1_IVG0
array 0 1 184 0 0 -415
timestamp 1704392934
transform 1 0 736 0 -1 498
box -17 -17 17 17
use via_M1_M2_0  MP1_IVS0
array 0 2 184 0 0 -415
timestamp 1704392934
transform 1 0 644 0 -1 747
box -17 -17 17 17
use via_M2_M3_0  NoName_0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704386899
transform 1 0 184 0 1 332
box -32 -17 32 17
use via_M2_M3_0  NoName_2
timestamp 1704386899
transform 1 0 184 0 1 498
box -32 -17 32 17
use via_M2_M3_0  NoName_3
timestamp 1704386899
transform 1 0 920 0 1 249
box -32 -17 32 17
use via_M2_M3_0  NoName_5
timestamp 1704386899
transform 1 0 920 0 1 581
box -32 -17 32 17
use via_M2_M3_0  NoName_6
timestamp 1704386899
transform 1 0 1012 0 1 332
box -32 -17 32 17
use via_M2_M3_0  NoName_10
timestamp 1704386899
transform 1 0 828 0 1 498
box -32 -17 32 17
use via_M1_M2_0  NoName_13
timestamp 1704392934
transform 1 0 552 0 1 581
box -17 -17 17 17
use via_M1_M2_0  NoName_15
timestamp 1704392934
transform 1 0 552 0 1 747
box -17 -17 17 17
use via_M1_M2_0  NoName_18
timestamp 1704392934
transform 1 0 552 0 1 249
box -17 -17 17 17
use via_M1_M2_0  NoName_20
timestamp 1704392934
transform 1 0 552 0 1 83
box -17 -17 17 17
<< labels >>
flabel metal1 1012 415 1012 415 0 FreeSans 512 90 0 0 EN
port 1 nsew
flabel metal1 828 415 828 415 0 FreeSans 512 90 0 0 ENB
port 2 nsew
flabel metal1 184 415 184 415 0 FreeSans 512 90 0 0 I
port 3 nsew
flabel metal1 920 415 920 415 0 FreeSans 512 90 0 0 O
port 4 nsew
flabel metal1 552 830 552 830 0 FreeSans 416 0 0 0 VDD
port 5 nsew
flabel metal1 552 0 552 0 0 FreeSans 416 0 0 0 VSS
port 6 nsew
<< end >>
