magic
tech sky130A
magscale 1 2
timestamp 1704394705
<< checkpaint >>
rect -1260 2116 2072 2156
rect -1294 -799 2072 2116
rect -1294 -1286 2030 -799
rect -1260 -1344 1996 -1286
<< locali >>
rect 66 713 118 864
rect 250 713 302 864
rect 434 713 486 864
rect 618 713 670 864
rect 139 564 597 598
rect 75 481 597 515
rect 75 315 597 349
rect 139 232 597 266
rect 66 -34 118 117
rect 250 -34 302 117
rect 434 -34 486 117
rect 618 -34 670 117
<< metal1 >>
rect 60 306 124 524
rect 152 223 216 607
rect 336 223 400 607
rect 520 223 584 607
<< metal2 >>
rect -34 804 770 856
rect -34 -26 770 26
use nmos130_fast_boundary  MN0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363493
transform 1 0 0 0 1 0
box 0 -84 92 280
use nmos130_fast_boundary  MN0_IBNDR0
timestamp 1704363493
transform 1 0 644 0 1 0
box 0 -84 92 280
use nmos130_fast_center_nf2  MN0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 2 184 0 0 415
timestamp 1704390143
transform 1 0 92 0 1 0
box -31 -84 215 362
use via_M1_M2_0  MN0_IVD0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 2 184 0 0 415
timestamp 1704392934
transform 1 0 184 0 1 249
box -17 -17 17 17
use via_M1_M2_0  MN0_IVG0
array 0 2 184 0 0 415
timestamp 1704392934
transform 1 0 184 0 1 332
box -17 -17 17 17
use via_M2_M3_M4  MN0_IVTIED0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 3 184 0 0 415
timestamp 1704389274
transform 1 0 92 0 1 0
box -32 -26 32 26
use pmos130_fast_boundary  MP0_IBNDL0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704363574
transform 1 0 0 0 -1 830
box 0 -66 168 369
use pmos130_fast_boundary  MP0_IBNDR0
timestamp 1704363574
transform 1 0 644 0 -1 830
box 0 -66 168 369
use pmos130_fast_center_nf2  MP0_IM0 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 2 184 0 0 -415
timestamp 1704364343
transform 1 0 92 0 -1 830
box -31 -66 215 369
use via_M1_M2_0  MP0_IVD0
array 0 2 184 0 0 -415
timestamp 1704392934
transform 1 0 184 0 -1 581
box -17 -17 17 17
use via_M1_M2_0  MP0_IVG0
array 0 2 184 0 0 -415
timestamp 1704392934
transform 1 0 184 0 -1 498
box -17 -17 17 17
use via_M2_M3_M4  MP0_IVTIED0
array 0 3 184 0 0 -415
timestamp 1704389274
transform 1 0 92 0 -1 830
box -32 -26 32 26
use via_M2_M3_0  NoName_1 /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1704386899
transform 1 0 92 0 1 332
box -32 -17 32 17
use via_M2_M3_0  NoName_3
timestamp 1704386899
transform 1 0 92 0 1 498
box -32 -17 32 17
use via_M2_M3_0  NoName_5
timestamp 1704386899
transform 1 0 184 0 1 249
box -32 -17 32 17
use via_M2_M3_0  NoName_7
timestamp 1704386899
transform 1 0 184 0 1 581
box -32 -17 32 17
use via_M2_M3_0  NoName_8
timestamp 1704386899
transform 1 0 368 0 1 249
box -32 -17 32 17
use via_M2_M3_0  NoName_10
timestamp 1704386899
transform 1 0 368 0 1 581
box -32 -17 32 17
use via_M2_M3_0  NoName_11
timestamp 1704386899
transform 1 0 552 0 1 249
box -32 -17 32 17
use via_M2_M3_0  NoName_13
timestamp 1704386899
transform 1 0 552 0 1 581
box -32 -17 32 17
<< labels >>
flabel metal1 92 415 92 415 0 FreeSans 512 90 0 0 I
port 1 nsew
flabel metal1 184 415 184 415 0 FreeSans 512 90 0 0 O:
port 2 nsew
flabel metal1 368 415 368 415 0 FreeSans 512 90 0 0 O:
port 3 nsew
flabel metal1 552 415 552 415 0 FreeSans 512 90 0 0 O:
port 4 nsew
flabel metal2 368 830 368 830 0 FreeSans 416 0 0 0 VDD
port 5 nsew
flabel metal2 368 0 368 0 0 FreeSans 416 0 0 0 VSS
port 6 nsew
<< end >>
