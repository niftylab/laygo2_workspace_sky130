magic
tech sky130A
timestamp 1704363523
<< pwell >>
rect 0 -42 92 140
<< properties >>
string FIXED_BBOX 0 0 92 207
<< end >>
