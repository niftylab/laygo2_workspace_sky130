magic
tech sky130A
magscale 1 2
timestamp 1679624521
<< checkpaint >>
rect -1300 -1325 2452 3337
<< metal2 >>
rect -40 1956 1192 2076
rect 258 978 750 1038
rect -40 -60 1192 60
<< metal3 >>
rect 114 720 174 1296
rect 834 432 894 1584
use logic_generated_inv_2x  inv0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/logic_generated
timestamp 1679560816
transform 1 0 0 0 1 0
box -40 -60 616 2076
use logic_generated_inv_2x  inv1
timestamp 1679560816
transform 1 0 576 0 1 0
box -40 -60 616 2076
use via_M2_M3_0  w1_net_w1_net_0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 288 0 1 1008
box -38 -38 38 38
use via_M2_M3_0  w1_net_w1_net_1
timestamp 1647525786
transform 1 0 720 0 1 1008
box -38 -38 38 38
<< labels >>
flabel metal3 144 1008 144 1008 0 FreeSans 480 90 0 0 I
port 1 nsew
flabel metal3 864 1008 864 1008 0 FreeSans 480 90 0 0 O
port 2 nsew
flabel metal2 576 2016 576 2016 0 FreeSans 960 0 0 0 VDD
port 3 nsew
flabel metal2 576 0 576 0 0 FreeSans 960 0 0 0 VSS
port 4 nsew
<< end >>
