magic
tech sky130A
magscale 1 2
timestamp 1679560830
<< checkpaint >>
rect -1300 3276 2432 3337
rect -1300 -268 2436 3276
rect -1300 -1325 2432 -268
<< metal1 >>
rect 114 1688 174 2056
rect 402 1688 462 2056
rect 690 1688 750 2056
rect 978 1688 1038 2056
rect 114 -40 174 328
rect 402 -40 462 328
rect 690 -40 750 328
rect 978 -40 1038 328
<< metal2 >>
rect -40 1956 1172 2076
rect 108 1554 468 1614
rect 720 1554 1008 1614
rect 108 1266 468 1326
rect 108 690 468 750
rect 108 402 468 462
rect 720 402 1008 462
rect -40 -60 1172 60
<< metal3 >>
rect 114 690 174 1326
use nmos13_fast_boundary  MN0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 144 1008
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 432 0 1 0
box 0 0 144 1008
use nmos13_fast_center_nf2  MN0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654175211
transform 1 0 144 0 1 0
box -92 286 380 756
use via_M1_M2_0  MN0_IVD0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 288 0 1 432
box -32 -32 32 32
use via_M1_M2_0  MN0_IVG0
timestamp 1647525606
transform 1 0 288 0 1 720
box -32 -32 32 32
use via_M1_M2_1  MN0_IVTIED0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 288 0 0 1008
timestamp 1647525606
transform 1 0 144 0 1 0
box -32 -32 32 32
use ntap_fast_boundary  MNT0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825115
transform 1 0 576 0 1 0
box 0 0 144 1024
use ntap_fast_boundary  MNT0_IBNDR0
timestamp 1655825115
transform 1 0 1008 0 1 0
box 0 0 144 1024
use ntap_fast_center_nf2_v2  MNT0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656694979
transform 1 0 720 0 1 0
box -72 286 360 684
use via_M1_M2_0  MNT0_IVTAP10
timestamp 1647525606
transform 1 0 864 0 1 432
box -32 -32 32 32
use via_M1_M2_1  MNT0_IVTIETAP10
array 0 1 288 0 0 1008
timestamp 1647525606
transform 1 0 720 0 1 0
box -32 -32 32 32
use pmos13_fast_boundary  MP0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 2016
box 0 0 144 1008
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 432 0 -1 2016
box 0 0 144 1008
use pmos13_fast_center_nf2  MP0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1654091791
transform 1 0 144 0 -1 2016
box -92 132 380 756
use via_M1_M2_0  MP0_IVD0
timestamp 1647525606
transform 1 0 288 0 -1 1584
box -32 -32 32 32
use via_M1_M2_0  MP0_IVG0
timestamp 1647525606
transform 1 0 288 0 -1 1296
box -32 -32 32 32
use via_M1_M2_1  MP0_IVTIED0
array 0 1 288 0 0 -1008
timestamp 1647525606
transform 1 0 144 0 -1 2016
box -32 -32 32 32
use ptap_fast_boundary  MPT0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825477
transform 1 0 576 0 -1 2016
box 0 0 168 1024
use ptap_fast_boundary  MPT0_IBNDR0
timestamp 1655825477
transform 1 0 1008 0 -1 2016
box 0 0 168 1024
use ptap_fast_center_nf2_v2  MPT0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656699071
transform 1 0 720 0 -1 2016
box -72 132 360 684
use via_M1_M2_0  MPT0_IVTAP10
timestamp 1647525606
transform 1 0 864 0 -1 1584
box -32 -32 32 32
use via_M1_M2_1  MPT0_IVTIETAP10
array 0 1 288 0 0 -1008
timestamp 1647525606
transform 1 0 720 0 -1 2016
box -32 -32 32 32
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 144 0 1 720
box -38 -38 38 38
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 144 0 1 1296
box -38 -38 38 38
<< labels >>
flabel metal3 144 1008 144 1008 0 FreeSans 480 90 0 0 I
port 1 nsew
flabel metal2 288 2016 288 2016 0 FreeSans 960 0 0 0 VDD
port 2 nsew
flabel metal2 288 0 288 0 0 FreeSans 960 0 0 0 VSS
port 3 nsew
<< end >>
