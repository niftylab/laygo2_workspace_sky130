magic
tech sky130A
timestamp 1679560818
<< checkpaint >>
rect -650 -660 3386 1668
<< metal1 >>
rect 57 844 87 1028
rect 201 844 231 1028
rect 345 844 375 1028
rect 489 844 519 1028
rect 633 844 663 1028
rect 777 844 807 1028
rect 921 844 951 1028
rect 1065 844 1095 1028
rect 1209 844 1239 1028
rect 1353 844 1383 1028
rect 1497 844 1527 1028
rect 1641 844 1671 1028
rect 1785 844 1815 1028
rect 1929 844 1959 1028
rect 2073 844 2103 1028
rect 2217 844 2247 1028
rect 2361 844 2391 1028
rect 2505 844 2535 1028
rect 2649 844 2679 1028
rect 57 -20 87 164
rect 201 -20 231 164
rect 345 -20 375 164
rect 489 -20 519 164
rect 633 -20 663 164
rect 777 -20 807 164
rect 921 -20 951 164
rect 1065 -20 1095 164
rect 1209 -20 1239 164
rect 1353 -20 1383 164
rect 1497 -20 1527 164
rect 1641 -20 1671 164
rect 1785 -20 1815 164
rect 1929 -20 1959 164
rect 2073 -20 2103 164
rect 2217 -20 2247 164
rect 2361 -20 2391 164
rect 2505 -20 2535 164
rect 2649 -20 2679 164
<< metal2 >>
rect -20 978 2756 1038
rect 106 777 2630 807
rect 62 633 2630 663
rect 62 345 2630 375
rect 106 201 2630 231
rect -20 -30 2756 30
<< metal3 >>
rect 57 345 87 663
rect 129 201 159 807
rect 273 201 303 807
rect 417 201 447 807
rect 561 201 591 807
rect 705 201 735 807
rect 849 201 879 807
rect 993 201 1023 807
rect 1137 201 1167 807
rect 1281 201 1311 807
rect 1425 201 1455 807
rect 1569 201 1599 807
rect 1713 201 1743 807
rect 1857 201 1887 807
rect 2001 201 2031 807
rect 2145 201 2175 807
rect 2289 201 2319 807
rect 2433 201 2463 807
rect 2577 201 2607 807
use nmos13_fast_boundary  MN0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 2664 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 17 144 0 0 504
timestamp 1654175211
transform 1 0 72 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN0_IVD0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 17 144 0 0 504
timestamp 1647525606
transform 1 0 144 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN0_IVG0
array 0 17 144 0 0 504
timestamp 1647525606
transform 1 0 144 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN0_IVTIED0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 18 144 0 0 504
timestamp 1647525606
transform 1 0 72 0 1 0
box -16 -16 16 16
use pmos13_fast_boundary  MP0_IBNDL0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 2664 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP0_IM0 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 17 144 0 0 -504
timestamp 1654091791
transform 1 0 72 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP0_IVD0
array 0 17 144 0 0 -504
timestamp 1647525606
transform 1 0 144 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP0_IVG0
array 0 17 144 0 0 -504
timestamp 1647525606
transform 1 0 144 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP0_IVTIED0
array 0 18 144 0 0 -504
timestamp 1647525606
transform 1 0 72 0 -1 1008
box -16 -16 16 16
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 72 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 72 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 144 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 144 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_8
timestamp 1647525786
transform 1 0 288 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_10
timestamp 1647525786
transform 1 0 288 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_11
timestamp 1647525786
transform 1 0 432 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_13
timestamp 1647525786
transform 1 0 432 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_14
timestamp 1647525786
transform 1 0 576 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_16
timestamp 1647525786
transform 1 0 576 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_17
timestamp 1647525786
transform 1 0 720 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_19
timestamp 1647525786
transform 1 0 720 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_20
timestamp 1647525786
transform 1 0 864 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_22
timestamp 1647525786
transform 1 0 864 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_23
timestamp 1647525786
transform 1 0 1008 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_25
timestamp 1647525786
transform 1 0 1008 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_26
timestamp 1647525786
transform 1 0 1152 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_28
timestamp 1647525786
transform 1 0 1152 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_29
timestamp 1647525786
transform 1 0 1296 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_31
timestamp 1647525786
transform 1 0 1296 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_32
timestamp 1647525786
transform 1 0 1440 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_34
timestamp 1647525786
transform 1 0 1440 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_35
timestamp 1647525786
transform 1 0 1584 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_37
timestamp 1647525786
transform 1 0 1584 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_38
timestamp 1647525786
transform 1 0 1728 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_40
timestamp 1647525786
transform 1 0 1728 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_41
timestamp 1647525786
transform 1 0 1872 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_43
timestamp 1647525786
transform 1 0 1872 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_44
timestamp 1647525786
transform 1 0 2016 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_46
timestamp 1647525786
transform 1 0 2016 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_47
timestamp 1647525786
transform 1 0 2160 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_49
timestamp 1647525786
transform 1 0 2160 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_50
timestamp 1647525786
transform 1 0 2304 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_52
timestamp 1647525786
transform 1 0 2304 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_53
timestamp 1647525786
transform 1 0 2448 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_55
timestamp 1647525786
transform 1 0 2448 0 1 792
box -19 -19 19 19
use via_M2_M3_0  NoName_56
timestamp 1647525786
transform 1 0 2592 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_58
timestamp 1647525786
transform 1 0 2592 0 1 792
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 I
port 24 nsew
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 O
port 25 nsew
flabel metal3 288 504 288 504 0 FreeSans 240 90 0 0 O
port 26 nsew
flabel metal3 432 504 432 504 0 FreeSans 240 90 0 0 O
port 27 nsew
flabel metal3 576 504 576 504 0 FreeSans 240 90 0 0 O
port 28 nsew
flabel metal3 720 504 720 504 0 FreeSans 240 90 0 0 O
port 29 nsew
flabel metal3 864 504 864 504 0 FreeSans 240 90 0 0 O
port 30 nsew
flabel metal3 1008 504 1008 504 0 FreeSans 240 90 0 0 O
port 31 nsew
flabel metal3 1152 504 1152 504 0 FreeSans 240 90 0 0 O
port 32 nsew
flabel metal3 1296 504 1296 504 0 FreeSans 240 90 0 0 O
port 33 nsew
flabel metal3 1728 504 1728 504 0 FreeSans 240 90 0 0 O
port 34 nsew
flabel metal3 2304 504 2304 504 0 FreeSans 240 90 0 0 O
port 35 nsew
flabel metal3 2592 504 2592 504 0 FreeSans 240 90 0 0 O
port 36 nsew
flabel metal3 144 504 144 504 0 FreeSans 240 90 0 0 O:
port 110 nsew
flabel metal3 288 504 288 504 0 FreeSans 240 90 0 0 O:
port 111 nsew
flabel metal3 432 504 432 504 0 FreeSans 240 90 0 0 O:
port 112 nsew
flabel metal3 576 504 576 504 0 FreeSans 240 90 0 0 O:
port 113 nsew
flabel metal3 720 504 720 504 0 FreeSans 240 90 0 0 O:
port 114 nsew
flabel metal3 864 504 864 504 0 FreeSans 240 90 0 0 O:
port 115 nsew
flabel metal3 1008 504 1008 504 0 FreeSans 240 90 0 0 O:
port 116 nsew
flabel metal3 1152 504 1152 504 0 FreeSans 240 90 0 0 O:
port 117 nsew
flabel metal3 1296 504 1296 504 0 FreeSans 240 90 0 0 O:
port 118 nsew
flabel metal3 1440 504 1440 504 0 FreeSans 240 90 0 0 O:
port 119 nsew
flabel metal3 1584 504 1584 504 0 FreeSans 240 90 0 0 O:
port 120 nsew
flabel metal3 1728 504 1728 504 0 FreeSans 240 90 0 0 O:
port 121 nsew
flabel metal3 1872 504 1872 504 0 FreeSans 240 90 0 0 O:
port 122 nsew
flabel metal3 2016 504 2016 504 0 FreeSans 240 90 0 0 O:
port 123 nsew
flabel metal3 2160 504 2160 504 0 FreeSans 240 90 0 0 O:
port 124 nsew
flabel metal3 2304 504 2304 504 0 FreeSans 240 90 0 0 O:
port 125 nsew
flabel metal3 2448 504 2448 504 0 FreeSans 240 90 0 0 O:
port 126 nsew
flabel metal3 2592 504 2592 504 0 FreeSans 240 90 0 0 O:
port 127 nsew
flabel metal2 144 1008 144 1008 0 FreeSans 480 0 0 0 VDD
port 140 nsew
flabel metal2 216 1008 216 1008 0 FreeSans 480 0 0 0 VDD
port 141 nsew
flabel metal2 288 1008 288 1008 0 FreeSans 480 0 0 0 VDD
port 142 nsew
flabel metal2 360 1008 360 1008 0 FreeSans 480 0 0 0 VDD
port 143 nsew
flabel metal2 432 1008 432 1008 0 FreeSans 480 0 0 0 VDD
port 144 nsew
flabel metal2 504 1008 504 1008 0 FreeSans 480 0 0 0 VDD
port 145 nsew
flabel metal2 576 1008 576 1008 0 FreeSans 480 0 0 0 VDD
port 146 nsew
flabel metal2 648 1008 648 1008 0 FreeSans 480 0 0 0 VDD
port 147 nsew
flabel metal2 720 1008 720 1008 0 FreeSans 480 0 0 0 VDD
port 148 nsew
flabel metal2 936 1008 936 1008 0 FreeSans 480 0 0 0 VDD
port 149 nsew
flabel metal2 1224 1008 1224 1008 0 FreeSans 480 0 0 0 VDD
port 150 nsew
flabel metal2 1368 1008 1368 1008 0 FreeSans 480 0 0 0 VDD
port 151 nsew
flabel metal2 144 0 144 0 0 FreeSans 480 0 0 0 VSS
port 164 nsew
flabel metal2 216 0 216 0 0 FreeSans 480 0 0 0 VSS
port 165 nsew
flabel metal2 288 0 288 0 0 FreeSans 480 0 0 0 VSS
port 166 nsew
flabel metal2 360 0 360 0 0 FreeSans 480 0 0 0 VSS
port 167 nsew
flabel metal2 432 0 432 0 0 FreeSans 480 0 0 0 VSS
port 168 nsew
flabel metal2 504 0 504 0 0 FreeSans 480 0 0 0 VSS
port 169 nsew
flabel metal2 576 0 576 0 0 FreeSans 480 0 0 0 VSS
port 170 nsew
flabel metal2 648 0 648 0 0 FreeSans 480 0 0 0 VSS
port 171 nsew
flabel metal2 720 0 720 0 0 FreeSans 480 0 0 0 VSS
port 172 nsew
flabel metal2 936 0 936 0 0 FreeSans 480 0 0 0 VSS
port 173 nsew
flabel metal2 1224 0 1224 0 0 FreeSans 480 0 0 0 VSS
port 174 nsew
flabel metal2 1368 0 1368 0 0 FreeSans 480 0 0 0 VSS
port 175 nsew
<< end >>
