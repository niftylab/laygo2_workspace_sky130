magic
tech sky130A
timestamp 1704389274
<< locali >>
rect -16 8 16 13
rect -16 -9 -9 8
rect 8 -9 16 8
rect -16 -13 16 -9
<< viali >>
rect -9 -9 8 8
<< metal1 >>
rect -16 -13 -13 13
rect 13 -13 16 13
<< via1 >>
rect -13 8 13 13
rect -13 -9 -9 8
rect -9 -9 8 8
rect 8 -9 13 8
rect -13 -13 13 -9
<< metal2 >>
rect -16 -13 -13 13
rect 13 -13 16 13
<< labels >>
flabel metal2 -13 -13 13 13 0 FreeSans 40 0 0 0 m2m1li
<< end >>
