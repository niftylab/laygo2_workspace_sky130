* SPICE3 file created from /WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense/nmos13_fast_center_nf2.ext - technology: sky130A

.subckt x/WORK/hjpark/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense/nmos13_fast_center_nf2
+ D0 G0 S0 S1 BODY
X0 D0 G0 S0 BODY sky130_fd_pr__nfet_01v8_lvt ad=2.394e+11p pd=1.98e+06u as=2.394e+11p ps=1.98e+06u w=420000u l=150000u
X1 D0 G0 S1 BODY sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.394e+11p ps=1.98e+06u w=420000u l=150000u
.ends

