magic
tech sky130A
timestamp 1679560847
<< checkpaint >>
rect -650 -660 2090 1668
<< metal2 >>
rect -20 978 1460 1038
rect 561 489 807 519
rect -20 -30 1460 30
<< metal3 >>
rect 57 360 87 648
rect 561 201 591 519
rect 777 345 807 519
rect 1281 216 1311 792
use logic_generated_inv_8x  inv0 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 0 0 1 0
box -20 -30 740 1038
use logic_generated_inv_8x  inv1
timestamp 1679560816
transform 1 0 720 0 1 0
box -20 -30 740 1038
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 576 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 792 0 1 504
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 I
port 1 nsew
flabel metal3 1296 504 1296 504 0 FreeSans 240 90 0 0 O
port 2 nsew
flabel metal2 720 1008 720 1008 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal2 720 0 720 0 0 FreeSans 480 0 0 0 VSS
port 4 nsew
<< end >>
