magic
tech sky130A
magscale 1 2
timestamp 1662802026
<< nwell >>
rect -92 132 380 684
<< pmos >>
rect 56 168 86 648
rect 200 168 230 648
<< pdiff >>
rect -56 578 56 648
rect -56 538 -20 578
rect 20 538 56 578
rect -56 478 56 538
rect -56 438 -20 478
rect 20 438 56 478
rect -56 378 56 438
rect -56 338 -20 378
rect 20 338 56 378
rect -56 278 56 338
rect -56 238 -20 278
rect 20 238 56 278
rect -56 168 56 238
rect 86 578 200 648
rect 86 538 124 578
rect 164 538 200 578
rect 86 478 200 538
rect 86 438 124 478
rect 164 438 200 478
rect 86 378 200 438
rect 86 338 124 378
rect 164 338 200 378
rect 86 278 200 338
rect 86 238 124 278
rect 164 238 200 278
rect 86 168 200 238
rect 230 578 344 648
rect 230 538 268 578
rect 308 538 344 578
rect 230 478 344 538
rect 230 438 268 478
rect 308 438 344 478
rect 230 378 344 438
rect 230 338 268 378
rect 308 338 344 378
rect 230 278 344 338
rect 230 238 268 278
rect 308 238 344 278
rect 230 168 344 238
<< pdiffc >>
rect -20 538 20 578
rect -20 438 20 478
rect -20 338 20 378
rect -20 238 20 278
rect 124 538 164 578
rect 124 438 164 478
rect 124 338 164 378
rect 124 238 164 278
rect 268 538 308 578
rect 268 438 308 478
rect 268 338 308 378
rect 268 238 308 278
<< poly >>
rect 56 737 230 756
rect 56 703 76 737
rect 110 703 184 737
rect 218 703 230 737
rect 56 684 230 703
rect 56 648 86 684
rect 200 648 230 684
rect 56 132 86 168
rect 200 132 230 168
<< polycont >>
rect 76 703 110 737
rect 184 703 218 737
<< locali >>
rect 56 737 230 756
rect 56 703 76 737
rect 110 703 184 737
rect 218 703 230 737
rect 56 684 230 703
rect -30 578 30 594
rect -30 538 -20 578
rect 20 538 30 578
rect -30 478 30 538
rect -30 438 -20 478
rect 20 438 30 478
rect -30 378 30 438
rect -30 338 -20 378
rect 20 338 30 378
rect -30 278 30 338
rect -30 238 -20 278
rect 20 238 30 278
rect -30 222 30 238
rect 114 578 174 594
rect 114 538 124 578
rect 164 538 174 578
rect 114 478 174 538
rect 114 438 124 478
rect 164 438 174 478
rect 114 378 174 438
rect 114 338 124 378
rect 164 338 174 378
rect 114 278 174 338
rect 114 238 124 278
rect 164 238 174 278
rect 114 222 174 238
rect 258 578 318 594
rect 258 538 268 578
rect 308 538 318 578
rect 258 478 318 538
rect 258 438 268 478
rect 308 438 318 478
rect 258 378 318 438
rect 258 338 268 378
rect 308 338 318 378
rect 258 278 318 338
rect 258 238 268 278
rect 308 238 318 278
rect 258 222 318 238
<< labels >>
flabel nwell -20 654 4 670 0 FreeSans 80 0 0 0 BODY
port 5 nsew
<< end >>
