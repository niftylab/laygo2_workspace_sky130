magic
tech sky130A
magscale 1 2
timestamp 1704386899
<< checkpaint >>
rect -1292 -1286 1292 1286
<< error_p >>
rect -17 -17 17 17
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -32 -17 -17 17
rect 17 -17 32 17
<< end >>
