magic
tech sky130A
timestamp 1679560857
<< checkpaint >>
rect -650 -660 3530 1668
<< metal2 >>
rect -20 978 2900 1038
rect 1281 489 1527 519
rect -20 -30 2900 30
<< metal3 >>
rect 57 360 87 648
rect 1281 201 1311 519
rect 1497 345 1527 519
rect 2721 216 2751 792
use logic_generated_inv_18x  inv0 magic_layout/logic_generated
timestamp 1679560816
transform 1 0 0 0 1 0
box -20 -30 1460 1038
use logic_generated_inv_18x  inv1
timestamp 1679560816
transform 1 0 1440 0 1 0
box -20 -30 1460 1038
use via_M2_M3_0  NoName_1 ~/WORK/sylee/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 1296 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 1512 0 1 504
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 I
port 1 nsew
flabel metal3 2736 504 2736 504 0 FreeSans 240 90 0 0 O
port 2 nsew
flabel metal2 1440 1008 1440 1008 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal2 1440 0 1440 0 0 FreeSans 480 0 0 0 VSS
port 4 nsew
<< end >>
