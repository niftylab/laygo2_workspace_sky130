magic
tech sky130A
timestamp 1704387567
<< labels >>
flabel space -13 -13 13 13 0 FreeSans 56 0 0 0 short
<< end >>
