magic
tech sky130A
timestamp 1655971500
<< checkpaint >>
rect -650 -660 4970 1668
<< metal2 >>
rect -20 978 4340 1038
rect -20 -30 4340 30
<< metal3 >>
rect 273 129 303 231
rect 489 129 519 375
rect 705 57 735 231
rect 1497 57 1527 375
rect 1569 129 1599 231
rect 1641 129 1671 375
rect 1785 273 1815 375
rect 1857 129 1887 375
rect 1929 129 1959 231
rect 2001 57 2031 375
rect 2217 201 2247 375
rect 2433 201 2463 303
rect 2721 273 2751 375
rect 3225 129 3255 375
rect 3297 129 3327 231
rect 3369 57 3399 375
rect 3513 273 3543 375
rect 3585 57 3615 375
rect 3657 129 3687 231
rect 3729 129 3759 375
rect 3945 201 3975 375
rect 4161 201 4191 303
<< metal4 >>
rect 1785 273 2751 303
rect 3513 273 4191 303
rect 1569 201 2247 231
rect 3297 201 3975 231
rect 273 129 3759 159
rect 705 57 3615 87
use via_M3_M4_0  NoName_1 skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 720 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_3
timestamp 1647526059
transform 1 0 1512 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_5
timestamp 1647526059
transform 1 0 3384 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_7
timestamp 1647526059
transform 1 0 2016 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_9
timestamp 1647526059
transform 1 0 3600 0 1 72
box -19 -19 19 19
use via_M3_M4_0  NoName_12
timestamp 1647526059
transform 1 0 288 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_14
timestamp 1647526059
transform 1 0 504 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_16
timestamp 1647526059
transform 1 0 1656 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_18
timestamp 1647526059
transform 1 0 3240 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_20
timestamp 1647526059
transform 1 0 1872 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_22
timestamp 1647526059
transform 1 0 3744 0 1 144
box -19 -19 19 19
use via_M3_M4_0  NoName_25
timestamp 1647526059
transform 1 0 2232 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_27
timestamp 1647526059
transform 1 0 1584 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_29
timestamp 1647526059
transform 1 0 1944 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_32
timestamp 1647526059
transform 1 0 3960 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_34
timestamp 1647526059
transform 1 0 3312 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_36
timestamp 1647526059
transform 1 0 3672 0 1 216
box -19 -19 19 19
use via_M3_M4_0  NoName_39
timestamp 1647526059
transform 1 0 2448 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_41
timestamp 1647526059
transform 1 0 2736 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_43
timestamp 1647526059
transform 1 0 1800 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_46
timestamp 1647526059
transform 1 0 4176 0 1 288
box -19 -19 19 19
use via_M3_M4_0  NoName_48
timestamp 1647526059
transform 1 0 3528 0 1 288
box -19 -19 19 19
use logic_generated_inv_4x  inv0
timestamp 1655971085
transform 1 0 0 0 1 0
box -20 -30 452 1038
use logic_generated_inv_4x  inv1
timestamp 1655971085
transform 1 0 432 0 1 0
box -20 -30 452 1038
use logic_generated_inv_4x  inv2
timestamp 1655971085
transform 1 0 2160 0 1 0
box -20 -30 452 1038
use logic_generated_inv_4x  inv3
timestamp 1655971085
transform 1 0 3888 0 1 0
box -20 -30 452 1038
use logic_generated_tinv_4x  tinv0
timestamp 1655971092
transform 1 0 864 0 1 0
box -20 -30 884 1038
use logic_generated_tinv_4x  tinv1
timestamp 1655971092
transform 1 0 2592 0 1 0
box -20 -30 884 1038
use logic_generated_tinv_small_1x  tinv_small0
timestamp 1655971095
transform 1 0 1728 0 1 0
box -20 -30 452 1038
use logic_generated_tinv_small_1x  tinv_small1
timestamp 1655971095
transform 1 0 3456 0 1 0
box -20 -30 452 1038
<< labels >>
flabel metal3 1008 504 1008 504 0 FreeSans 240 90 0 0 I
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 CLK
flabel metal3 4176 504 4176 504 0 FreeSans 240 90 0 0 O
flabel metal2 2160 0 2160 0 0 FreeSans 480 0 0 0 VSS
flabel metal2 2160 1008 2160 1008 0 FreeSans 480 0 0 0 VDD
<< end >>
