magic
tech sky130A
timestamp 1654176054
<< pwell >>
rect -46 186 190 342
<< nmoslvt >>
rect 28 204 43 324
rect 100 204 115 324
<< ndiff >>
rect -28 299 28 324
rect -28 279 -10 299
rect 10 279 28 299
rect -28 249 28 279
rect -28 229 -10 249
rect 10 229 28 249
rect -28 204 28 229
rect 43 299 100 324
rect 43 279 62 299
rect 82 279 100 299
rect 43 249 100 279
rect 43 229 62 249
rect 82 229 100 249
rect 43 204 100 229
rect 115 299 172 324
rect 115 279 134 299
rect 154 279 172 299
rect 115 249 172 279
rect 115 229 134 249
rect 154 229 172 249
rect 115 204 172 229
<< ndiffc >>
rect -10 279 10 299
rect -10 229 10 249
rect 62 279 82 299
rect 62 229 82 249
rect 134 279 154 299
rect 134 229 154 249
<< poly >>
rect -17 369 43 378
rect -17 351 -6 369
rect 12 351 43 369
rect -17 342 43 351
rect 28 324 43 342
rect 100 369 160 378
rect 100 351 133 369
rect 151 351 160 369
rect 100 342 160 351
rect 100 324 115 342
rect 28 186 43 204
rect 100 186 115 204
<< polycont >>
rect -6 351 12 369
rect 133 351 151 369
<< locali >>
rect -17 369 28 378
rect -17 351 -6 369
rect 12 351 28 369
rect -17 342 28 351
rect 115 369 160 378
rect 115 351 133 369
rect 151 351 160 369
rect 115 342 160 351
rect -15 299 15 307
rect -15 279 -10 299
rect 10 279 15 299
rect -15 249 15 279
rect -15 229 -10 249
rect 10 229 15 249
rect -15 221 15 229
rect 57 299 87 307
rect 57 279 62 299
rect 82 279 87 299
rect 57 249 87 279
rect 57 229 62 249
rect 82 229 87 249
rect 57 221 87 229
rect 129 299 159 307
rect 129 279 134 299
rect 154 279 159 299
rect 129 249 159 279
rect 129 229 134 249
rect 154 229 159 249
rect 129 221 159 229
<< viali >>
rect -6 351 12 369
rect 133 351 151 369
rect -10 279 10 299
rect -10 229 10 249
rect 62 279 82 299
rect 62 229 82 249
rect 134 279 154 299
rect 134 229 154 249
<< metal1 >>
rect -17 369 28 378
rect -17 351 -6 369
rect 12 351 28 369
rect -17 342 28 351
rect 115 369 160 378
rect 115 351 133 369
rect 151 351 160 369
rect 115 342 160 351
rect -15 299 15 307
rect -15 279 -10 299
rect 10 279 15 299
rect -15 249 15 279
rect -15 229 -10 249
rect 10 229 15 249
rect -15 144 15 229
rect 57 299 87 307
rect 57 279 62 299
rect 82 279 87 299
rect 57 249 87 279
rect 57 229 62 249
rect 82 229 87 249
rect 57 221 87 229
rect 129 299 159 307
rect 129 279 134 299
rect 154 279 159 299
rect 129 249 159 279
rect 129 229 134 249
rect 154 229 159 249
rect 129 144 159 229
<< labels >>
flabel metal1 -17 342 28 378 0 FreeSans 80 0 0 0 G0
port 2 nsew
flabel metal1 115 342 160 378 0 FreeSans 80 0 0 0 G1
port 3 nsew
flabel metal1 -15 144 15 307 0 FreeSans 80 0 0 0 S0
port 4 nsew
rlabel pwell -20 327 -5 338 1 BODY
port 6 nsew
flabel metal1 129 144 159 307 0 FreeSans 80 0 0 0 D0
port 1 e
<< end >>
